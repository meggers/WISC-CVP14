module picker();
  
endmodule
