module CVP14(output [15:0] Addr, output RD, output WR, output V, output U, output [15:0] dataOut, 
             input Reset, input Clk1, input Clk2, input [15:0] DataIn);
            
VectorRegFile vrf();
ScalarRegFile srf();
ALU alu();

endmodule
