
module CVP14 ( Addr, RD, WR, V, dataOut, Reset, Clk1, Clk2, DataIn );
  output [15:0] Addr;
  output [15:0] dataOut;
  input [15:0] DataIn;
  input Reset, Clk1, Clk2;
  output RD, WR, V;
  wire   N152, N153, N155, overflow, N1457, N1458, N1459, N1460, N1461, N1462,
         N1463, N1464, N1465, N1466, N1467, N1468, N1469, N1470, N1471, N1472,
         N1473, N1474, N1475, N1476, N1477, N1478, N1479, N1480, N1481, N1482,
         N1483, N1810, N1811, N1812, N1813, N1814, N1815, N1816, N1817, N1818,
         N1819, N1820, N1821, N1822, N1823, N1824, N1825, N4133, N4134, N4135,
         N4136, N4137, N4138, N4139, N4140, N4141, N4142, N4143, N4144, N4145,
         N4146, N4147, N4148, N4149, N4153, N4154, N4155, N4156, N4157, N4158,
         N4159, N4160, N4161, N4162, N4163, N4164, N4165, N4166, N4167, N4168,
         N4169, N4170, N4171, N4172, N4173, N4174, N4175, N4176, N4177, N4178,
         N4179, N4180, N4181, N4182, N4183, N4184, N4185, N4186, N4187, N4188,
         N4189, N4190, N4191, N4192, N4193, N4194, N4195, N4196, N4197, N4198,
         N4199, N4200, N4201, N4202, N4203, N4204, N4205, N4206, N4207, N4208,
         N4209, N4210, N4211, N4212, N4213, N4214, N4215, N4216, N4217, N4218,
         N4219, N4220, N4221, N4222, N4223, N4224, N4225, N4226, N4227, N4228,
         N4229, N4230, N4231, N4233, N4234, N4235, N4236, N4237, N4238, N4239,
         N4240, N4241, N4242, N4243, N4244, N4245, N4246, N4247, N4248, N4249,
         N4250, N4251, N4252, N4253, N4254, N4255, N4256, N4257, N4258, N4259,
         N4260, N4261, N4262, N4263, N4264, N4265, N4266, N4267, N4268, N4269,
         N4270, N4271, N4272, N4273, N4274, N4275, N4276, N4277, N4278, N4279,
         N4280, N4281, N4282, N4283, N4284, N4285, N4286, N4287, N4288, N4289,
         N4290, N4291, N4292, N4293, N4294, N4295, N4296, N4297, N4298, N4299,
         N4300, N4301, N4302, N4303, N4304, N4305, N4306, N4307, N4308, N4309,
         N4310, N4311, N4312, N4313, N4314, N4315, N4316, N4317, N4318, N4319,
         N4320, N4321, N4322, N4323, N4324, N4325, N4326, N4327, N4328, N4329,
         N4330, N4331, N4333, N4334, N4335, N4336, N4337, N4338, N4339, N4340,
         N4341, N4342, N4343, N4344, N4345, N4346, N4347, N4348, N4349, N4350,
         N4351, N4352, N4353, N4354, N4355, N4356, N4357, N4358, N4359, N4360,
         N4361, N4362, N4363, N4364, N4365, N4366, N4367, N4368, N4369, N4370,
         N4371, N4372, N4373, N4374, N4375, N4376, N4377, N4378, N4379, N4380,
         N4381, N4382, N4383, N4384, N4385, N4386, N4387, N4388, N4389, N4390,
         N4391, N4392, N4393, N4394, N4395, N4396, N4397, N4398, N4399, N4400,
         N4401, N4402, N4403, N4404, N4405, N4406, N4407, N4408, N4409, N4410,
         N4411, N4412, N4413, N4414, N4415, N4416, N4417, N4418, N4419, N4420,
         N4421, N4422, N4423, N4424, N4425, N4426, N4427, N4428, N4429, N4430,
         N4431, N4433, N4434, N4435, N4436, N4437, N4438, N4439, N4440, N4441,
         N4442, N4443, N4444, N4445, N4446, N4447, N4448, N4449, N4450, N4451,
         N4452, N4453, N4454, N4455, N4456, N4457, N4458, N4459, N4460, N4461,
         N4462, N4463, N4464, N4465, N4466, N4467, N4468, N4469, N4470, N4471,
         N4472, N4473, N4474, \vrf/N296 , \vrf/N293 , \vrf/N290 , \vrf/N287 ,
         \vrf/N284 , \vrf/N281 , \vrf/N278 , \vrf/N275 , \vrf/N274 ,
         \vrf/N273 , \vrf/N272 , \vrf/N271 , \vrf/N270 , \vrf/N269 ,
         \vrf/N268 , \vrf/N267 , \vrf/N266 , \vrf/N265 , \vrf/N264 ,
         \vrf/N263 , \vrf/N262 , \vrf/N261 , \vrf/N260 , \vrf/N259 ,
         \vrf/N258 , \vrf/N257 , \vrf/N256 , \vrf/N255 , \vrf/N254 ,
         \vrf/N253 , \vrf/N252 , \vrf/N251 , \vrf/N250 , \vrf/N249 ,
         \vrf/N248 , \vrf/N247 , \vrf/N246 , \vrf/N245 , \vrf/N244 ,
         \vrf/N243 , \vrf/N242 , \vrf/N241 , \vrf/N240 , \vrf/N239 ,
         \vrf/N238 , \vrf/N237 , \vrf/N236 , \vrf/N235 , \vrf/N234 ,
         \vrf/N233 , \vrf/N232 , \vrf/N231 , \vrf/N230 , \vrf/N229 ,
         \vrf/N228 , \vrf/N227 , \vrf/N226 , \vrf/N225 , \vrf/N224 ,
         \vrf/N223 , \vrf/N222 , \vrf/N221 , \vrf/N220 , \vrf/N219 ,
         \vrf/N218 , \vrf/N217 , \vrf/N216 , \vrf/N215 , \vrf/N214 ,
         \vrf/N213 , \vrf/N212 , \vrf/N211 , \vrf/N210 , \vrf/N209 ,
         \vrf/N208 , \vrf/N207 , \vrf/N206 , \vrf/N205 , \vrf/N204 ,
         \vrf/N203 , \vrf/N202 , \vrf/N201 , \vrf/N200 , \vrf/N199 ,
         \vrf/N198 , \vrf/N197 , \vrf/N196 , \vrf/N195 , \vrf/N194 ,
         \vrf/N193 , \vrf/N192 , \vrf/N191 , \vrf/N190 , \vrf/N189 ,
         \vrf/N188 , \vrf/N187 , \vrf/N186 , \vrf/N185 , \vrf/N184 ,
         \vrf/N183 , \vrf/N182 , \vrf/N181 , \vrf/N180 , \vrf/N179 ,
         \vrf/N178 , \vrf/N177 , \vrf/N176 , \vrf/N175 , \vrf/N174 ,
         \vrf/N173 , \vrf/N172 , \vrf/N171 , \vrf/N170 , \vrf/N169 ,
         \vrf/N168 , \vrf/N167 , \vrf/N166 , \vrf/N165 , \vrf/N164 ,
         \vrf/N163 , \vrf/N162 , \vrf/N161 , \vrf/N160 , \vrf/N159 ,
         \vrf/N158 , \vrf/N157 , \vrf/N156 , \vrf/N155 , \vrf/N154 ,
         \vrf/N153 , \vrf/N152 , \vrf/N151 , \vrf/N150 , \vrf/N149 ,
         \vrf/N148 , \vrf/N147 , \vrf/N146 , \vrf/N145 , \vrf/N144 ,
         \vrf/N143 , \vrf/N142 , \vrf/N141 , \vrf/N140 , \vrf/N139 ,
         \vrf/N138 , \vrf/N137 , \vrf/N136 , \vrf/N135 , \vrf/N134 ,
         \vrf/N133 , \vrf/N132 , \vrf/N131 , \vrf/N130 , \vrf/N129 ,
         \vrf/N128 , \vrf/N127 , \vrf/N126 , \vrf/N125 , \vrf/N124 ,
         \vrf/N123 , \vrf/N122 , \vrf/N121 , \vrf/N120 , \vrf/N119 ,
         \vrf/N118 , \vrf/N116 , \vrf/N115 , \vrf/N114 , \vrf/N113 ,
         \vrf/N112 , \vrf/N111 , \vrf/N110 , \vrf/N109 , \vrf/N108 ,
         \vrf/N107 , \vrf/N106 , \vrf/N105 , \vrf/N104 , \vrf/N103 ,
         \vrf/N102 , \vrf/N101 , \vrf/N100 , \vrf/N99 , \vrf/N98 , \vrf/N97 ,
         \vrf/N96 , \vrf/N95 , \vrf/N94 , \vrf/N93 , \vrf/N92 , \vrf/N91 ,
         \vrf/N90 , \vrf/N89 , \vrf/N88 , \vrf/N87 , \vrf/N86 , \vrf/N85 ,
         \vrf/N84 , \vrf/N83 , \vrf/N82 , \vrf/N81 , \vrf/N80 , \vrf/N79 ,
         \vrf/N78 , \vrf/N77 , \vrf/N76 , \vrf/N75 , \vrf/N74 , \vrf/N73 ,
         \vrf/N72 , \vrf/N71 , \vrf/N70 , \vrf/N69 , \vrf/N68 , \vrf/N67 ,
         \vrf/N66 , \vrf/N65 , \vrf/N64 , \vrf/N63 , \vrf/N62 , \vrf/N61 ,
         \vrf/N60 , \vrf/N59 , \vrf/N58 , \vrf/N57 , \vrf/N56 , \vrf/N55 ,
         \vrf/N54 , \vrf/N53 , \vrf/N52 , \vrf/N51 , \vrf/N50 , \vrf/N49 ,
         \vrf/N48 , \vrf/N47 , \vrf/N46 , \vrf/N45 , \vrf/N44 , \vrf/N43 ,
         \vrf/N42 , \vrf/N41 , \vrf/N40 , \vrf/N39 , \vrf/N38 , \vrf/N37 ,
         \vrf/N36 , \vrf/N35 , \vrf/N34 , \vrf/N33 , \vrf/N32 , \vrf/N31 ,
         \vrf/N30 , \vrf/N29 , \vrf/N28 , \vrf/N27 , \vrf/N26 , \vrf/N25 ,
         \vrf/N24 , \vrf/N23 , \vrf/N22 , \vrf/N21 , \vrf/N20 , \vrf/N19 ,
         \vrf/N18 , \vrf/regTable[7][0] , \vrf/regTable[7][1] ,
         \vrf/regTable[7][2] , \vrf/regTable[7][3] , \vrf/regTable[7][4] ,
         \vrf/regTable[7][5] , \vrf/regTable[7][6] , \vrf/regTable[7][7] ,
         \vrf/regTable[7][8] , \vrf/regTable[7][9] , \vrf/regTable[7][10] ,
         \vrf/regTable[7][11] , \vrf/regTable[7][12] , \vrf/regTable[7][13] ,
         \vrf/regTable[7][14] , \vrf/regTable[7][15] , \vrf/regTable[7][16] ,
         \vrf/regTable[7][17] , \vrf/regTable[7][18] , \vrf/regTable[7][19] ,
         \vrf/regTable[7][20] , \vrf/regTable[7][21] , \vrf/regTable[7][22] ,
         \vrf/regTable[7][23] , \vrf/regTable[7][24] , \vrf/regTable[7][25] ,
         \vrf/regTable[7][26] , \vrf/regTable[7][27] , \vrf/regTable[7][28] ,
         \vrf/regTable[7][29] , \vrf/regTable[7][30] , \vrf/regTable[7][31] ,
         \vrf/regTable[7][32] , \vrf/regTable[7][33] , \vrf/regTable[7][34] ,
         \vrf/regTable[7][35] , \vrf/regTable[7][36] , \vrf/regTable[7][37] ,
         \vrf/regTable[7][38] , \vrf/regTable[7][39] , \vrf/regTable[7][40] ,
         \vrf/regTable[7][41] , \vrf/regTable[7][42] , \vrf/regTable[7][43] ,
         \vrf/regTable[7][44] , \vrf/regTable[7][45] , \vrf/regTable[7][46] ,
         \vrf/regTable[7][47] , \vrf/regTable[7][48] , \vrf/regTable[7][49] ,
         \vrf/regTable[7][50] , \vrf/regTable[7][51] , \vrf/regTable[7][52] ,
         \vrf/regTable[7][53] , \vrf/regTable[7][54] , \vrf/regTable[7][55] ,
         \vrf/regTable[7][56] , \vrf/regTable[7][57] , \vrf/regTable[7][58] ,
         \vrf/regTable[7][59] , \vrf/regTable[7][60] , \vrf/regTable[7][61] ,
         \vrf/regTable[7][62] , \vrf/regTable[7][63] , \vrf/regTable[7][64] ,
         \vrf/regTable[7][65] , \vrf/regTable[7][66] , \vrf/regTable[7][67] ,
         \vrf/regTable[7][68] , \vrf/regTable[7][69] , \vrf/regTable[7][70] ,
         \vrf/regTable[7][71] , \vrf/regTable[7][72] , \vrf/regTable[7][73] ,
         \vrf/regTable[7][74] , \vrf/regTable[7][75] , \vrf/regTable[7][76] ,
         \vrf/regTable[7][77] , \vrf/regTable[7][78] , \vrf/regTable[7][79] ,
         \vrf/regTable[7][80] , \vrf/regTable[7][81] , \vrf/regTable[7][82] ,
         \vrf/regTable[7][83] , \vrf/regTable[7][84] , \vrf/regTable[7][85] ,
         \vrf/regTable[7][86] , \vrf/regTable[7][87] , \vrf/regTable[7][88] ,
         \vrf/regTable[7][89] , \vrf/regTable[7][90] , \vrf/regTable[7][91] ,
         \vrf/regTable[7][92] , \vrf/regTable[7][93] , \vrf/regTable[7][94] ,
         \vrf/regTable[7][95] , \vrf/regTable[7][96] , \vrf/regTable[7][97] ,
         \vrf/regTable[7][98] , \vrf/regTable[7][99] , \vrf/regTable[7][100] ,
         \vrf/regTable[7][101] , \vrf/regTable[7][102] ,
         \vrf/regTable[7][103] , \vrf/regTable[7][104] ,
         \vrf/regTable[7][105] , \vrf/regTable[7][106] ,
         \vrf/regTable[7][107] , \vrf/regTable[7][108] ,
         \vrf/regTable[7][109] , \vrf/regTable[7][110] ,
         \vrf/regTable[7][111] , \vrf/regTable[7][112] ,
         \vrf/regTable[7][113] , \vrf/regTable[7][114] ,
         \vrf/regTable[7][115] , \vrf/regTable[7][116] ,
         \vrf/regTable[7][117] , \vrf/regTable[7][118] ,
         \vrf/regTable[7][119] , \vrf/regTable[7][120] ,
         \vrf/regTable[7][121] , \vrf/regTable[7][122] ,
         \vrf/regTable[7][123] , \vrf/regTable[7][124] ,
         \vrf/regTable[7][125] , \vrf/regTable[7][126] ,
         \vrf/regTable[7][127] , \vrf/regTable[7][128] ,
         \vrf/regTable[7][129] , \vrf/regTable[7][130] ,
         \vrf/regTable[7][131] , \vrf/regTable[7][132] ,
         \vrf/regTable[7][133] , \vrf/regTable[7][134] ,
         \vrf/regTable[7][135] , \vrf/regTable[7][136] ,
         \vrf/regTable[7][137] , \vrf/regTable[7][138] ,
         \vrf/regTable[7][139] , \vrf/regTable[7][140] ,
         \vrf/regTable[7][141] , \vrf/regTable[7][142] ,
         \vrf/regTable[7][143] , \vrf/regTable[7][144] ,
         \vrf/regTable[7][145] , \vrf/regTable[7][146] ,
         \vrf/regTable[7][147] , \vrf/regTable[7][148] ,
         \vrf/regTable[7][149] , \vrf/regTable[7][150] ,
         \vrf/regTable[7][151] , \vrf/regTable[7][152] ,
         \vrf/regTable[7][153] , \vrf/regTable[7][154] ,
         \vrf/regTable[7][155] , \vrf/regTable[7][156] ,
         \vrf/regTable[7][157] , \vrf/regTable[7][158] ,
         \vrf/regTable[7][159] , \vrf/regTable[7][160] ,
         \vrf/regTable[7][161] , \vrf/regTable[7][162] ,
         \vrf/regTable[7][163] , \vrf/regTable[7][164] ,
         \vrf/regTable[7][165] , \vrf/regTable[7][166] ,
         \vrf/regTable[7][167] , \vrf/regTable[7][168] ,
         \vrf/regTable[7][169] , \vrf/regTable[7][170] ,
         \vrf/regTable[7][171] , \vrf/regTable[7][172] ,
         \vrf/regTable[7][173] , \vrf/regTable[7][174] ,
         \vrf/regTable[7][175] , \vrf/regTable[7][176] ,
         \vrf/regTable[7][177] , \vrf/regTable[7][178] ,
         \vrf/regTable[7][179] , \vrf/regTable[7][180] ,
         \vrf/regTable[7][181] , \vrf/regTable[7][182] ,
         \vrf/regTable[7][183] , \vrf/regTable[7][184] ,
         \vrf/regTable[7][185] , \vrf/regTable[7][186] ,
         \vrf/regTable[7][187] , \vrf/regTable[7][188] ,
         \vrf/regTable[7][189] , \vrf/regTable[7][190] ,
         \vrf/regTable[7][191] , \vrf/regTable[7][192] ,
         \vrf/regTable[7][193] , \vrf/regTable[7][194] ,
         \vrf/regTable[7][195] , \vrf/regTable[7][196] ,
         \vrf/regTable[7][197] , \vrf/regTable[7][198] ,
         \vrf/regTable[7][199] , \vrf/regTable[7][200] ,
         \vrf/regTable[7][201] , \vrf/regTable[7][202] ,
         \vrf/regTable[7][203] , \vrf/regTable[7][204] ,
         \vrf/regTable[7][205] , \vrf/regTable[7][206] ,
         \vrf/regTable[7][207] , \vrf/regTable[7][208] ,
         \vrf/regTable[7][209] , \vrf/regTable[7][210] ,
         \vrf/regTable[7][211] , \vrf/regTable[7][212] ,
         \vrf/regTable[7][213] , \vrf/regTable[7][214] ,
         \vrf/regTable[7][215] , \vrf/regTable[7][216] ,
         \vrf/regTable[7][217] , \vrf/regTable[7][218] ,
         \vrf/regTable[7][219] , \vrf/regTable[7][220] ,
         \vrf/regTable[7][221] , \vrf/regTable[7][222] ,
         \vrf/regTable[7][223] , \vrf/regTable[7][224] ,
         \vrf/regTable[7][225] , \vrf/regTable[7][226] ,
         \vrf/regTable[7][227] , \vrf/regTable[7][228] ,
         \vrf/regTable[7][229] , \vrf/regTable[7][230] ,
         \vrf/regTable[7][231] , \vrf/regTable[7][232] ,
         \vrf/regTable[7][233] , \vrf/regTable[7][234] ,
         \vrf/regTable[7][235] , \vrf/regTable[7][236] ,
         \vrf/regTable[7][237] , \vrf/regTable[7][238] ,
         \vrf/regTable[7][239] , \vrf/regTable[7][240] ,
         \vrf/regTable[7][241] , \vrf/regTable[7][242] ,
         \vrf/regTable[7][243] , \vrf/regTable[7][244] ,
         \vrf/regTable[7][245] , \vrf/regTable[7][246] ,
         \vrf/regTable[7][247] , \vrf/regTable[7][248] ,
         \vrf/regTable[7][249] , \vrf/regTable[7][250] ,
         \vrf/regTable[7][251] , \vrf/regTable[7][252] ,
         \vrf/regTable[7][253] , \vrf/regTable[7][254] ,
         \vrf/regTable[7][255] , \vrf/regTable[6][0] , \vrf/regTable[6][1] ,
         \vrf/regTable[6][2] , \vrf/regTable[6][3] , \vrf/regTable[6][4] ,
         \vrf/regTable[6][5] , \vrf/regTable[6][6] , \vrf/regTable[6][7] ,
         \vrf/regTable[6][8] , \vrf/regTable[6][9] , \vrf/regTable[6][10] ,
         \vrf/regTable[6][11] , \vrf/regTable[6][12] , \vrf/regTable[6][13] ,
         \vrf/regTable[6][14] , \vrf/regTable[6][15] , \vrf/regTable[6][16] ,
         \vrf/regTable[6][17] , \vrf/regTable[6][18] , \vrf/regTable[6][19] ,
         \vrf/regTable[6][20] , \vrf/regTable[6][21] , \vrf/regTable[6][22] ,
         \vrf/regTable[6][23] , \vrf/regTable[6][24] , \vrf/regTable[6][25] ,
         \vrf/regTable[6][26] , \vrf/regTable[6][27] , \vrf/regTable[6][28] ,
         \vrf/regTable[6][29] , \vrf/regTable[6][30] , \vrf/regTable[6][31] ,
         \vrf/regTable[6][32] , \vrf/regTable[6][33] , \vrf/regTable[6][34] ,
         \vrf/regTable[6][35] , \vrf/regTable[6][36] , \vrf/regTable[6][37] ,
         \vrf/regTable[6][38] , \vrf/regTable[6][39] , \vrf/regTable[6][40] ,
         \vrf/regTable[6][41] , \vrf/regTable[6][42] , \vrf/regTable[6][43] ,
         \vrf/regTable[6][44] , \vrf/regTable[6][45] , \vrf/regTable[6][46] ,
         \vrf/regTable[6][47] , \vrf/regTable[6][48] , \vrf/regTable[6][49] ,
         \vrf/regTable[6][50] , \vrf/regTable[6][51] , \vrf/regTable[6][52] ,
         \vrf/regTable[6][53] , \vrf/regTable[6][54] , \vrf/regTable[6][55] ,
         \vrf/regTable[6][56] , \vrf/regTable[6][57] , \vrf/regTable[6][58] ,
         \vrf/regTable[6][59] , \vrf/regTable[6][60] , \vrf/regTable[6][61] ,
         \vrf/regTable[6][62] , \vrf/regTable[6][63] , \vrf/regTable[6][64] ,
         \vrf/regTable[6][65] , \vrf/regTable[6][66] , \vrf/regTable[6][67] ,
         \vrf/regTable[6][68] , \vrf/regTable[6][69] , \vrf/regTable[6][70] ,
         \vrf/regTable[6][71] , \vrf/regTable[6][72] , \vrf/regTable[6][73] ,
         \vrf/regTable[6][74] , \vrf/regTable[6][75] , \vrf/regTable[6][76] ,
         \vrf/regTable[6][77] , \vrf/regTable[6][78] , \vrf/regTable[6][79] ,
         \vrf/regTable[6][80] , \vrf/regTable[6][81] , \vrf/regTable[6][82] ,
         \vrf/regTable[6][83] , \vrf/regTable[6][84] , \vrf/regTable[6][85] ,
         \vrf/regTable[6][86] , \vrf/regTable[6][87] , \vrf/regTable[6][88] ,
         \vrf/regTable[6][89] , \vrf/regTable[6][90] , \vrf/regTable[6][91] ,
         \vrf/regTable[6][92] , \vrf/regTable[6][93] , \vrf/regTable[6][94] ,
         \vrf/regTable[6][95] , \vrf/regTable[6][96] , \vrf/regTable[6][97] ,
         \vrf/regTable[6][98] , \vrf/regTable[6][99] , \vrf/regTable[6][100] ,
         \vrf/regTable[6][101] , \vrf/regTable[6][102] ,
         \vrf/regTable[6][103] , \vrf/regTable[6][104] ,
         \vrf/regTable[6][105] , \vrf/regTable[6][106] ,
         \vrf/regTable[6][107] , \vrf/regTable[6][108] ,
         \vrf/regTable[6][109] , \vrf/regTable[6][110] ,
         \vrf/regTable[6][111] , \vrf/regTable[6][112] ,
         \vrf/regTable[6][113] , \vrf/regTable[6][114] ,
         \vrf/regTable[6][115] , \vrf/regTable[6][116] ,
         \vrf/regTable[6][117] , \vrf/regTable[6][118] ,
         \vrf/regTable[6][119] , \vrf/regTable[6][120] ,
         \vrf/regTable[6][121] , \vrf/regTable[6][122] ,
         \vrf/regTable[6][123] , \vrf/regTable[6][124] ,
         \vrf/regTable[6][125] , \vrf/regTable[6][126] ,
         \vrf/regTable[6][127] , \vrf/regTable[6][128] ,
         \vrf/regTable[6][129] , \vrf/regTable[6][130] ,
         \vrf/regTable[6][131] , \vrf/regTable[6][132] ,
         \vrf/regTable[6][133] , \vrf/regTable[6][134] ,
         \vrf/regTable[6][135] , \vrf/regTable[6][136] ,
         \vrf/regTable[6][137] , \vrf/regTable[6][138] ,
         \vrf/regTable[6][139] , \vrf/regTable[6][140] ,
         \vrf/regTable[6][141] , \vrf/regTable[6][142] ,
         \vrf/regTable[6][143] , \vrf/regTable[6][144] ,
         \vrf/regTable[6][145] , \vrf/regTable[6][146] ,
         \vrf/regTable[6][147] , \vrf/regTable[6][148] ,
         \vrf/regTable[6][149] , \vrf/regTable[6][150] ,
         \vrf/regTable[6][151] , \vrf/regTable[6][152] ,
         \vrf/regTable[6][153] , \vrf/regTable[6][154] ,
         \vrf/regTable[6][155] , \vrf/regTable[6][156] ,
         \vrf/regTable[6][157] , \vrf/regTable[6][158] ,
         \vrf/regTable[6][159] , \vrf/regTable[6][160] ,
         \vrf/regTable[6][161] , \vrf/regTable[6][162] ,
         \vrf/regTable[6][163] , \vrf/regTable[6][164] ,
         \vrf/regTable[6][165] , \vrf/regTable[6][166] ,
         \vrf/regTable[6][167] , \vrf/regTable[6][168] ,
         \vrf/regTable[6][169] , \vrf/regTable[6][170] ,
         \vrf/regTable[6][171] , \vrf/regTable[6][172] ,
         \vrf/regTable[6][173] , \vrf/regTable[6][174] ,
         \vrf/regTable[6][175] , \vrf/regTable[6][176] ,
         \vrf/regTable[6][177] , \vrf/regTable[6][178] ,
         \vrf/regTable[6][179] , \vrf/regTable[6][180] ,
         \vrf/regTable[6][181] , \vrf/regTable[6][182] ,
         \vrf/regTable[6][183] , \vrf/regTable[6][184] ,
         \vrf/regTable[6][185] , \vrf/regTable[6][186] ,
         \vrf/regTable[6][187] , \vrf/regTable[6][188] ,
         \vrf/regTable[6][189] , \vrf/regTable[6][190] ,
         \vrf/regTable[6][191] , \vrf/regTable[6][192] ,
         \vrf/regTable[6][193] , \vrf/regTable[6][194] ,
         \vrf/regTable[6][195] , \vrf/regTable[6][196] ,
         \vrf/regTable[6][197] , \vrf/regTable[6][198] ,
         \vrf/regTable[6][199] , \vrf/regTable[6][200] ,
         \vrf/regTable[6][201] , \vrf/regTable[6][202] ,
         \vrf/regTable[6][203] , \vrf/regTable[6][204] ,
         \vrf/regTable[6][205] , \vrf/regTable[6][206] ,
         \vrf/regTable[6][207] , \vrf/regTable[6][208] ,
         \vrf/regTable[6][209] , \vrf/regTable[6][210] ,
         \vrf/regTable[6][211] , \vrf/regTable[6][212] ,
         \vrf/regTable[6][213] , \vrf/regTable[6][214] ,
         \vrf/regTable[6][215] , \vrf/regTable[6][216] ,
         \vrf/regTable[6][217] , \vrf/regTable[6][218] ,
         \vrf/regTable[6][219] , \vrf/regTable[6][220] ,
         \vrf/regTable[6][221] , \vrf/regTable[6][222] ,
         \vrf/regTable[6][223] , \vrf/regTable[6][224] ,
         \vrf/regTable[6][225] , \vrf/regTable[6][226] ,
         \vrf/regTable[6][227] , \vrf/regTable[6][228] ,
         \vrf/regTable[6][229] , \vrf/regTable[6][230] ,
         \vrf/regTable[6][231] , \vrf/regTable[6][232] ,
         \vrf/regTable[6][233] , \vrf/regTable[6][234] ,
         \vrf/regTable[6][235] , \vrf/regTable[6][236] ,
         \vrf/regTable[6][237] , \vrf/regTable[6][238] ,
         \vrf/regTable[6][239] , \vrf/regTable[6][240] ,
         \vrf/regTable[6][241] , \vrf/regTable[6][242] ,
         \vrf/regTable[6][243] , \vrf/regTable[6][244] ,
         \vrf/regTable[6][245] , \vrf/regTable[6][246] ,
         \vrf/regTable[6][247] , \vrf/regTable[6][248] ,
         \vrf/regTable[6][249] , \vrf/regTable[6][250] ,
         \vrf/regTable[6][251] , \vrf/regTable[6][252] ,
         \vrf/regTable[6][253] , \vrf/regTable[6][254] ,
         \vrf/regTable[6][255] , \vrf/regTable[5][0] , \vrf/regTable[5][1] ,
         \vrf/regTable[5][2] , \vrf/regTable[5][3] , \vrf/regTable[5][4] ,
         \vrf/regTable[5][5] , \vrf/regTable[5][6] , \vrf/regTable[5][7] ,
         \vrf/regTable[5][8] , \vrf/regTable[5][9] , \vrf/regTable[5][10] ,
         \vrf/regTable[5][11] , \vrf/regTable[5][12] , \vrf/regTable[5][13] ,
         \vrf/regTable[5][14] , \vrf/regTable[5][15] , \vrf/regTable[5][16] ,
         \vrf/regTable[5][17] , \vrf/regTable[5][18] , \vrf/regTable[5][19] ,
         \vrf/regTable[5][20] , \vrf/regTable[5][21] , \vrf/regTable[5][22] ,
         \vrf/regTable[5][23] , \vrf/regTable[5][24] , \vrf/regTable[5][25] ,
         \vrf/regTable[5][26] , \vrf/regTable[5][27] , \vrf/regTable[5][28] ,
         \vrf/regTable[5][29] , \vrf/regTable[5][30] , \vrf/regTable[5][31] ,
         \vrf/regTable[5][32] , \vrf/regTable[5][33] , \vrf/regTable[5][34] ,
         \vrf/regTable[5][35] , \vrf/regTable[5][36] , \vrf/regTable[5][37] ,
         \vrf/regTable[5][38] , \vrf/regTable[5][39] , \vrf/regTable[5][40] ,
         \vrf/regTable[5][41] , \vrf/regTable[5][42] , \vrf/regTable[5][43] ,
         \vrf/regTable[5][44] , \vrf/regTable[5][45] , \vrf/regTable[5][46] ,
         \vrf/regTable[5][47] , \vrf/regTable[5][48] , \vrf/regTable[5][49] ,
         \vrf/regTable[5][50] , \vrf/regTable[5][51] , \vrf/regTable[5][52] ,
         \vrf/regTable[5][53] , \vrf/regTable[5][54] , \vrf/regTable[5][55] ,
         \vrf/regTable[5][56] , \vrf/regTable[5][57] , \vrf/regTable[5][58] ,
         \vrf/regTable[5][59] , \vrf/regTable[5][60] , \vrf/regTable[5][61] ,
         \vrf/regTable[5][62] , \vrf/regTable[5][63] , \vrf/regTable[5][64] ,
         \vrf/regTable[5][65] , \vrf/regTable[5][66] , \vrf/regTable[5][67] ,
         \vrf/regTable[5][68] , \vrf/regTable[5][69] , \vrf/regTable[5][70] ,
         \vrf/regTable[5][71] , \vrf/regTable[5][72] , \vrf/regTable[5][73] ,
         \vrf/regTable[5][74] , \vrf/regTable[5][75] , \vrf/regTable[5][76] ,
         \vrf/regTable[5][77] , \vrf/regTable[5][78] , \vrf/regTable[5][79] ,
         \vrf/regTable[5][80] , \vrf/regTable[5][81] , \vrf/regTable[5][82] ,
         \vrf/regTable[5][83] , \vrf/regTable[5][84] , \vrf/regTable[5][85] ,
         \vrf/regTable[5][86] , \vrf/regTable[5][87] , \vrf/regTable[5][88] ,
         \vrf/regTable[5][89] , \vrf/regTable[5][90] , \vrf/regTable[5][91] ,
         \vrf/regTable[5][92] , \vrf/regTable[5][93] , \vrf/regTable[5][94] ,
         \vrf/regTable[5][95] , \vrf/regTable[5][96] , \vrf/regTable[5][97] ,
         \vrf/regTable[5][98] , \vrf/regTable[5][99] , \vrf/regTable[5][100] ,
         \vrf/regTable[5][101] , \vrf/regTable[5][102] ,
         \vrf/regTable[5][103] , \vrf/regTable[5][104] ,
         \vrf/regTable[5][105] , \vrf/regTable[5][106] ,
         \vrf/regTable[5][107] , \vrf/regTable[5][108] ,
         \vrf/regTable[5][109] , \vrf/regTable[5][110] ,
         \vrf/regTable[5][111] , \vrf/regTable[5][112] ,
         \vrf/regTable[5][113] , \vrf/regTable[5][114] ,
         \vrf/regTable[5][115] , \vrf/regTable[5][116] ,
         \vrf/regTable[5][117] , \vrf/regTable[5][118] ,
         \vrf/regTable[5][119] , \vrf/regTable[5][120] ,
         \vrf/regTable[5][121] , \vrf/regTable[5][122] ,
         \vrf/regTable[5][123] , \vrf/regTable[5][124] ,
         \vrf/regTable[5][125] , \vrf/regTable[5][126] ,
         \vrf/regTable[5][127] , \vrf/regTable[5][128] ,
         \vrf/regTable[5][129] , \vrf/regTable[5][130] ,
         \vrf/regTable[5][131] , \vrf/regTable[5][132] ,
         \vrf/regTable[5][133] , \vrf/regTable[5][134] ,
         \vrf/regTable[5][135] , \vrf/regTable[5][136] ,
         \vrf/regTable[5][137] , \vrf/regTable[5][138] ,
         \vrf/regTable[5][139] , \vrf/regTable[5][140] ,
         \vrf/regTable[5][141] , \vrf/regTable[5][142] ,
         \vrf/regTable[5][143] , \vrf/regTable[5][144] ,
         \vrf/regTable[5][145] , \vrf/regTable[5][146] ,
         \vrf/regTable[5][147] , \vrf/regTable[5][148] ,
         \vrf/regTable[5][149] , \vrf/regTable[5][150] ,
         \vrf/regTable[5][151] , \vrf/regTable[5][152] ,
         \vrf/regTable[5][153] , \vrf/regTable[5][154] ,
         \vrf/regTable[5][155] , \vrf/regTable[5][156] ,
         \vrf/regTable[5][157] , \vrf/regTable[5][158] ,
         \vrf/regTable[5][159] , \vrf/regTable[5][160] ,
         \vrf/regTable[5][161] , \vrf/regTable[5][162] ,
         \vrf/regTable[5][163] , \vrf/regTable[5][164] ,
         \vrf/regTable[5][165] , \vrf/regTable[5][166] ,
         \vrf/regTable[5][167] , \vrf/regTable[5][168] ,
         \vrf/regTable[5][169] , \vrf/regTable[5][170] ,
         \vrf/regTable[5][171] , \vrf/regTable[5][172] ,
         \vrf/regTable[5][173] , \vrf/regTable[5][174] ,
         \vrf/regTable[5][175] , \vrf/regTable[5][176] ,
         \vrf/regTable[5][177] , \vrf/regTable[5][178] ,
         \vrf/regTable[5][179] , \vrf/regTable[5][180] ,
         \vrf/regTable[5][181] , \vrf/regTable[5][182] ,
         \vrf/regTable[5][183] , \vrf/regTable[5][184] ,
         \vrf/regTable[5][185] , \vrf/regTable[5][186] ,
         \vrf/regTable[5][187] , \vrf/regTable[5][188] ,
         \vrf/regTable[5][189] , \vrf/regTable[5][190] ,
         \vrf/regTable[5][191] , \vrf/regTable[5][192] ,
         \vrf/regTable[5][193] , \vrf/regTable[5][194] ,
         \vrf/regTable[5][195] , \vrf/regTable[5][196] ,
         \vrf/regTable[5][197] , \vrf/regTable[5][198] ,
         \vrf/regTable[5][199] , \vrf/regTable[5][200] ,
         \vrf/regTable[5][201] , \vrf/regTable[5][202] ,
         \vrf/regTable[5][203] , \vrf/regTable[5][204] ,
         \vrf/regTable[5][205] , \vrf/regTable[5][206] ,
         \vrf/regTable[5][207] , \vrf/regTable[5][208] ,
         \vrf/regTable[5][209] , \vrf/regTable[5][210] ,
         \vrf/regTable[5][211] , \vrf/regTable[5][212] ,
         \vrf/regTable[5][213] , \vrf/regTable[5][214] ,
         \vrf/regTable[5][215] , \vrf/regTable[5][216] ,
         \vrf/regTable[5][217] , \vrf/regTable[5][218] ,
         \vrf/regTable[5][219] , \vrf/regTable[5][220] ,
         \vrf/regTable[5][221] , \vrf/regTable[5][222] ,
         \vrf/regTable[5][223] , \vrf/regTable[5][224] ,
         \vrf/regTable[5][225] , \vrf/regTable[5][226] ,
         \vrf/regTable[5][227] , \vrf/regTable[5][228] ,
         \vrf/regTable[5][229] , \vrf/regTable[5][230] ,
         \vrf/regTable[5][231] , \vrf/regTable[5][232] ,
         \vrf/regTable[5][233] , \vrf/regTable[5][234] ,
         \vrf/regTable[5][235] , \vrf/regTable[5][236] ,
         \vrf/regTable[5][237] , \vrf/regTable[5][238] ,
         \vrf/regTable[5][239] , \vrf/regTable[5][240] ,
         \vrf/regTable[5][241] , \vrf/regTable[5][242] ,
         \vrf/regTable[5][243] , \vrf/regTable[5][244] ,
         \vrf/regTable[5][245] , \vrf/regTable[5][246] ,
         \vrf/regTable[5][247] , \vrf/regTable[5][248] ,
         \vrf/regTable[5][249] , \vrf/regTable[5][250] ,
         \vrf/regTable[5][251] , \vrf/regTable[5][252] ,
         \vrf/regTable[5][253] , \vrf/regTable[5][254] ,
         \vrf/regTable[5][255] , \vrf/regTable[4][0] , \vrf/regTable[4][1] ,
         \vrf/regTable[4][2] , \vrf/regTable[4][3] , \vrf/regTable[4][4] ,
         \vrf/regTable[4][5] , \vrf/regTable[4][6] , \vrf/regTable[4][7] ,
         \vrf/regTable[4][8] , \vrf/regTable[4][9] , \vrf/regTable[4][10] ,
         \vrf/regTable[4][11] , \vrf/regTable[4][12] , \vrf/regTable[4][13] ,
         \vrf/regTable[4][14] , \vrf/regTable[4][15] , \vrf/regTable[4][16] ,
         \vrf/regTable[4][17] , \vrf/regTable[4][18] , \vrf/regTable[4][19] ,
         \vrf/regTable[4][20] , \vrf/regTable[4][21] , \vrf/regTable[4][22] ,
         \vrf/regTable[4][23] , \vrf/regTable[4][24] , \vrf/regTable[4][25] ,
         \vrf/regTable[4][26] , \vrf/regTable[4][27] , \vrf/regTable[4][28] ,
         \vrf/regTable[4][29] , \vrf/regTable[4][30] , \vrf/regTable[4][31] ,
         \vrf/regTable[4][32] , \vrf/regTable[4][33] , \vrf/regTable[4][34] ,
         \vrf/regTable[4][35] , \vrf/regTable[4][36] , \vrf/regTable[4][37] ,
         \vrf/regTable[4][38] , \vrf/regTable[4][39] , \vrf/regTable[4][40] ,
         \vrf/regTable[4][41] , \vrf/regTable[4][42] , \vrf/regTable[4][43] ,
         \vrf/regTable[4][44] , \vrf/regTable[4][45] , \vrf/regTable[4][46] ,
         \vrf/regTable[4][47] , \vrf/regTable[4][48] , \vrf/regTable[4][49] ,
         \vrf/regTable[4][50] , \vrf/regTable[4][51] , \vrf/regTable[4][52] ,
         \vrf/regTable[4][53] , \vrf/regTable[4][54] , \vrf/regTable[4][55] ,
         \vrf/regTable[4][56] , \vrf/regTable[4][57] , \vrf/regTable[4][58] ,
         \vrf/regTable[4][59] , \vrf/regTable[4][60] , \vrf/regTable[4][61] ,
         \vrf/regTable[4][62] , \vrf/regTable[4][63] , \vrf/regTable[4][64] ,
         \vrf/regTable[4][65] , \vrf/regTable[4][66] , \vrf/regTable[4][67] ,
         \vrf/regTable[4][68] , \vrf/regTable[4][69] , \vrf/regTable[4][70] ,
         \vrf/regTable[4][71] , \vrf/regTable[4][72] , \vrf/regTable[4][73] ,
         \vrf/regTable[4][74] , \vrf/regTable[4][75] , \vrf/regTable[4][76] ,
         \vrf/regTable[4][77] , \vrf/regTable[4][78] , \vrf/regTable[4][79] ,
         \vrf/regTable[4][80] , \vrf/regTable[4][81] , \vrf/regTable[4][82] ,
         \vrf/regTable[4][83] , \vrf/regTable[4][84] , \vrf/regTable[4][85] ,
         \vrf/regTable[4][86] , \vrf/regTable[4][87] , \vrf/regTable[4][88] ,
         \vrf/regTable[4][89] , \vrf/regTable[4][90] , \vrf/regTable[4][91] ,
         \vrf/regTable[4][92] , \vrf/regTable[4][93] , \vrf/regTable[4][94] ,
         \vrf/regTable[4][95] , \vrf/regTable[4][96] , \vrf/regTable[4][97] ,
         \vrf/regTable[4][98] , \vrf/regTable[4][99] , \vrf/regTable[4][100] ,
         \vrf/regTable[4][101] , \vrf/regTable[4][102] ,
         \vrf/regTable[4][103] , \vrf/regTable[4][104] ,
         \vrf/regTable[4][105] , \vrf/regTable[4][106] ,
         \vrf/regTable[4][107] , \vrf/regTable[4][108] ,
         \vrf/regTable[4][109] , \vrf/regTable[4][110] ,
         \vrf/regTable[4][111] , \vrf/regTable[4][112] ,
         \vrf/regTable[4][113] , \vrf/regTable[4][114] ,
         \vrf/regTable[4][115] , \vrf/regTable[4][116] ,
         \vrf/regTable[4][117] , \vrf/regTable[4][118] ,
         \vrf/regTable[4][119] , \vrf/regTable[4][120] ,
         \vrf/regTable[4][121] , \vrf/regTable[4][122] ,
         \vrf/regTable[4][123] , \vrf/regTable[4][124] ,
         \vrf/regTable[4][125] , \vrf/regTable[4][126] ,
         \vrf/regTable[4][127] , \vrf/regTable[4][128] ,
         \vrf/regTable[4][129] , \vrf/regTable[4][130] ,
         \vrf/regTable[4][131] , \vrf/regTable[4][132] ,
         \vrf/regTable[4][133] , \vrf/regTable[4][134] ,
         \vrf/regTable[4][135] , \vrf/regTable[4][136] ,
         \vrf/regTable[4][137] , \vrf/regTable[4][138] ,
         \vrf/regTable[4][139] , \vrf/regTable[4][140] ,
         \vrf/regTable[4][141] , \vrf/regTable[4][142] ,
         \vrf/regTable[4][143] , \vrf/regTable[4][144] ,
         \vrf/regTable[4][145] , \vrf/regTable[4][146] ,
         \vrf/regTable[4][147] , \vrf/regTable[4][148] ,
         \vrf/regTable[4][149] , \vrf/regTable[4][150] ,
         \vrf/regTable[4][151] , \vrf/regTable[4][152] ,
         \vrf/regTable[4][153] , \vrf/regTable[4][154] ,
         \vrf/regTable[4][155] , \vrf/regTable[4][156] ,
         \vrf/regTable[4][157] , \vrf/regTable[4][158] ,
         \vrf/regTable[4][159] , \vrf/regTable[4][160] ,
         \vrf/regTable[4][161] , \vrf/regTable[4][162] ,
         \vrf/regTable[4][163] , \vrf/regTable[4][164] ,
         \vrf/regTable[4][165] , \vrf/regTable[4][166] ,
         \vrf/regTable[4][167] , \vrf/regTable[4][168] ,
         \vrf/regTable[4][169] , \vrf/regTable[4][170] ,
         \vrf/regTable[4][171] , \vrf/regTable[4][172] ,
         \vrf/regTable[4][173] , \vrf/regTable[4][174] ,
         \vrf/regTable[4][175] , \vrf/regTable[4][176] ,
         \vrf/regTable[4][177] , \vrf/regTable[4][178] ,
         \vrf/regTable[4][179] , \vrf/regTable[4][180] ,
         \vrf/regTable[4][181] , \vrf/regTable[4][182] ,
         \vrf/regTable[4][183] , \vrf/regTable[4][184] ,
         \vrf/regTable[4][185] , \vrf/regTable[4][186] ,
         \vrf/regTable[4][187] , \vrf/regTable[4][188] ,
         \vrf/regTable[4][189] , \vrf/regTable[4][190] ,
         \vrf/regTable[4][191] , \vrf/regTable[4][192] ,
         \vrf/regTable[4][193] , \vrf/regTable[4][194] ,
         \vrf/regTable[4][195] , \vrf/regTable[4][196] ,
         \vrf/regTable[4][197] , \vrf/regTable[4][198] ,
         \vrf/regTable[4][199] , \vrf/regTable[4][200] ,
         \vrf/regTable[4][201] , \vrf/regTable[4][202] ,
         \vrf/regTable[4][203] , \vrf/regTable[4][204] ,
         \vrf/regTable[4][205] , \vrf/regTable[4][206] ,
         \vrf/regTable[4][207] , \vrf/regTable[4][208] ,
         \vrf/regTable[4][209] , \vrf/regTable[4][210] ,
         \vrf/regTable[4][211] , \vrf/regTable[4][212] ,
         \vrf/regTable[4][213] , \vrf/regTable[4][214] ,
         \vrf/regTable[4][215] , \vrf/regTable[4][216] ,
         \vrf/regTable[4][217] , \vrf/regTable[4][218] ,
         \vrf/regTable[4][219] , \vrf/regTable[4][220] ,
         \vrf/regTable[4][221] , \vrf/regTable[4][222] ,
         \vrf/regTable[4][223] , \vrf/regTable[4][224] ,
         \vrf/regTable[4][225] , \vrf/regTable[4][226] ,
         \vrf/regTable[4][227] , \vrf/regTable[4][228] ,
         \vrf/regTable[4][229] , \vrf/regTable[4][230] ,
         \vrf/regTable[4][231] , \vrf/regTable[4][232] ,
         \vrf/regTable[4][233] , \vrf/regTable[4][234] ,
         \vrf/regTable[4][235] , \vrf/regTable[4][236] ,
         \vrf/regTable[4][237] , \vrf/regTable[4][238] ,
         \vrf/regTable[4][239] , \vrf/regTable[4][240] ,
         \vrf/regTable[4][241] , \vrf/regTable[4][242] ,
         \vrf/regTable[4][243] , \vrf/regTable[4][244] ,
         \vrf/regTable[4][245] , \vrf/regTable[4][246] ,
         \vrf/regTable[4][247] , \vrf/regTable[4][248] ,
         \vrf/regTable[4][249] , \vrf/regTable[4][250] ,
         \vrf/regTable[4][251] , \vrf/regTable[4][252] ,
         \vrf/regTable[4][253] , \vrf/regTable[4][254] ,
         \vrf/regTable[4][255] , \vrf/regTable[3][0] , \vrf/regTable[3][1] ,
         \vrf/regTable[3][2] , \vrf/regTable[3][3] , \vrf/regTable[3][4] ,
         \vrf/regTable[3][5] , \vrf/regTable[3][6] , \vrf/regTable[3][7] ,
         \vrf/regTable[3][8] , \vrf/regTable[3][9] , \vrf/regTable[3][10] ,
         \vrf/regTable[3][11] , \vrf/regTable[3][12] , \vrf/regTable[3][13] ,
         \vrf/regTable[3][14] , \vrf/regTable[3][15] , \vrf/regTable[3][16] ,
         \vrf/regTable[3][17] , \vrf/regTable[3][18] , \vrf/regTable[3][19] ,
         \vrf/regTable[3][20] , \vrf/regTable[3][21] , \vrf/regTable[3][22] ,
         \vrf/regTable[3][23] , \vrf/regTable[3][24] , \vrf/regTable[3][25] ,
         \vrf/regTable[3][26] , \vrf/regTable[3][27] , \vrf/regTable[3][28] ,
         \vrf/regTable[3][29] , \vrf/regTable[3][30] , \vrf/regTable[3][31] ,
         \vrf/regTable[3][32] , \vrf/regTable[3][33] , \vrf/regTable[3][34] ,
         \vrf/regTable[3][35] , \vrf/regTable[3][36] , \vrf/regTable[3][37] ,
         \vrf/regTable[3][38] , \vrf/regTable[3][39] , \vrf/regTable[3][40] ,
         \vrf/regTable[3][41] , \vrf/regTable[3][42] , \vrf/regTable[3][43] ,
         \vrf/regTable[3][44] , \vrf/regTable[3][45] , \vrf/regTable[3][46] ,
         \vrf/regTable[3][47] , \vrf/regTable[3][48] , \vrf/regTable[3][49] ,
         \vrf/regTable[3][50] , \vrf/regTable[3][51] , \vrf/regTable[3][52] ,
         \vrf/regTable[3][53] , \vrf/regTable[3][54] , \vrf/regTable[3][55] ,
         \vrf/regTable[3][56] , \vrf/regTable[3][57] , \vrf/regTable[3][58] ,
         \vrf/regTable[3][59] , \vrf/regTable[3][60] , \vrf/regTable[3][61] ,
         \vrf/regTable[3][62] , \vrf/regTable[3][63] , \vrf/regTable[3][64] ,
         \vrf/regTable[3][65] , \vrf/regTable[3][66] , \vrf/regTable[3][67] ,
         \vrf/regTable[3][68] , \vrf/regTable[3][69] , \vrf/regTable[3][70] ,
         \vrf/regTable[3][71] , \vrf/regTable[3][72] , \vrf/regTable[3][73] ,
         \vrf/regTable[3][74] , \vrf/regTable[3][75] , \vrf/regTable[3][76] ,
         \vrf/regTable[3][77] , \vrf/regTable[3][78] , \vrf/regTable[3][79] ,
         \vrf/regTable[3][80] , \vrf/regTable[3][81] , \vrf/regTable[3][82] ,
         \vrf/regTable[3][83] , \vrf/regTable[3][84] , \vrf/regTable[3][85] ,
         \vrf/regTable[3][86] , \vrf/regTable[3][87] , \vrf/regTable[3][88] ,
         \vrf/regTable[3][89] , \vrf/regTable[3][90] , \vrf/regTable[3][91] ,
         \vrf/regTable[3][92] , \vrf/regTable[3][93] , \vrf/regTable[3][94] ,
         \vrf/regTable[3][95] , \vrf/regTable[3][96] , \vrf/regTable[3][97] ,
         \vrf/regTable[3][98] , \vrf/regTable[3][99] , \vrf/regTable[3][100] ,
         \vrf/regTable[3][101] , \vrf/regTable[3][102] ,
         \vrf/regTable[3][103] , \vrf/regTable[3][104] ,
         \vrf/regTable[3][105] , \vrf/regTable[3][106] ,
         \vrf/regTable[3][107] , \vrf/regTable[3][108] ,
         \vrf/regTable[3][109] , \vrf/regTable[3][110] ,
         \vrf/regTable[3][111] , \vrf/regTable[3][112] ,
         \vrf/regTable[3][113] , \vrf/regTable[3][114] ,
         \vrf/regTable[3][115] , \vrf/regTable[3][116] ,
         \vrf/regTable[3][117] , \vrf/regTable[3][118] ,
         \vrf/regTable[3][119] , \vrf/regTable[3][120] ,
         \vrf/regTable[3][121] , \vrf/regTable[3][122] ,
         \vrf/regTable[3][123] , \vrf/regTable[3][124] ,
         \vrf/regTable[3][125] , \vrf/regTable[3][126] ,
         \vrf/regTable[3][127] , \vrf/regTable[3][128] ,
         \vrf/regTable[3][129] , \vrf/regTable[3][130] ,
         \vrf/regTable[3][131] , \vrf/regTable[3][132] ,
         \vrf/regTable[3][133] , \vrf/regTable[3][134] ,
         \vrf/regTable[3][135] , \vrf/regTable[3][136] ,
         \vrf/regTable[3][137] , \vrf/regTable[3][138] ,
         \vrf/regTable[3][139] , \vrf/regTable[3][140] ,
         \vrf/regTable[3][141] , \vrf/regTable[3][142] ,
         \vrf/regTable[3][143] , \vrf/regTable[3][144] ,
         \vrf/regTable[3][145] , \vrf/regTable[3][146] ,
         \vrf/regTable[3][147] , \vrf/regTable[3][148] ,
         \vrf/regTable[3][149] , \vrf/regTable[3][150] ,
         \vrf/regTable[3][151] , \vrf/regTable[3][152] ,
         \vrf/regTable[3][153] , \vrf/regTable[3][154] ,
         \vrf/regTable[3][155] , \vrf/regTable[3][156] ,
         \vrf/regTable[3][157] , \vrf/regTable[3][158] ,
         \vrf/regTable[3][159] , \vrf/regTable[3][160] ,
         \vrf/regTable[3][161] , \vrf/regTable[3][162] ,
         \vrf/regTable[3][163] , \vrf/regTable[3][164] ,
         \vrf/regTable[3][165] , \vrf/regTable[3][166] ,
         \vrf/regTable[3][167] , \vrf/regTable[3][168] ,
         \vrf/regTable[3][169] , \vrf/regTable[3][170] ,
         \vrf/regTable[3][171] , \vrf/regTable[3][172] ,
         \vrf/regTable[3][173] , \vrf/regTable[3][174] ,
         \vrf/regTable[3][175] , \vrf/regTable[3][176] ,
         \vrf/regTable[3][177] , \vrf/regTable[3][178] ,
         \vrf/regTable[3][179] , \vrf/regTable[3][180] ,
         \vrf/regTable[3][181] , \vrf/regTable[3][182] ,
         \vrf/regTable[3][183] , \vrf/regTable[3][184] ,
         \vrf/regTable[3][185] , \vrf/regTable[3][186] ,
         \vrf/regTable[3][187] , \vrf/regTable[3][188] ,
         \vrf/regTable[3][189] , \vrf/regTable[3][190] ,
         \vrf/regTable[3][191] , \vrf/regTable[3][192] ,
         \vrf/regTable[3][193] , \vrf/regTable[3][194] ,
         \vrf/regTable[3][195] , \vrf/regTable[3][196] ,
         \vrf/regTable[3][197] , \vrf/regTable[3][198] ,
         \vrf/regTable[3][199] , \vrf/regTable[3][200] ,
         \vrf/regTable[3][201] , \vrf/regTable[3][202] ,
         \vrf/regTable[3][203] , \vrf/regTable[3][204] ,
         \vrf/regTable[3][205] , \vrf/regTable[3][206] ,
         \vrf/regTable[3][207] , \vrf/regTable[3][208] ,
         \vrf/regTable[3][209] , \vrf/regTable[3][210] ,
         \vrf/regTable[3][211] , \vrf/regTable[3][212] ,
         \vrf/regTable[3][213] , \vrf/regTable[3][214] ,
         \vrf/regTable[3][215] , \vrf/regTable[3][216] ,
         \vrf/regTable[3][217] , \vrf/regTable[3][218] ,
         \vrf/regTable[3][219] , \vrf/regTable[3][220] ,
         \vrf/regTable[3][221] , \vrf/regTable[3][222] ,
         \vrf/regTable[3][223] , \vrf/regTable[3][224] ,
         \vrf/regTable[3][225] , \vrf/regTable[3][226] ,
         \vrf/regTable[3][227] , \vrf/regTable[3][228] ,
         \vrf/regTable[3][229] , \vrf/regTable[3][230] ,
         \vrf/regTable[3][231] , \vrf/regTable[3][232] ,
         \vrf/regTable[3][233] , \vrf/regTable[3][234] ,
         \vrf/regTable[3][235] , \vrf/regTable[3][236] ,
         \vrf/regTable[3][237] , \vrf/regTable[3][238] ,
         \vrf/regTable[3][239] , \vrf/regTable[3][240] ,
         \vrf/regTable[3][241] , \vrf/regTable[3][242] ,
         \vrf/regTable[3][243] , \vrf/regTable[3][244] ,
         \vrf/regTable[3][245] , \vrf/regTable[3][246] ,
         \vrf/regTable[3][247] , \vrf/regTable[3][248] ,
         \vrf/regTable[3][249] , \vrf/regTable[3][250] ,
         \vrf/regTable[3][251] , \vrf/regTable[3][252] ,
         \vrf/regTable[3][253] , \vrf/regTable[3][254] ,
         \vrf/regTable[3][255] , \vrf/regTable[2][0] , \vrf/regTable[2][1] ,
         \vrf/regTable[2][2] , \vrf/regTable[2][3] , \vrf/regTable[2][4] ,
         \vrf/regTable[2][5] , \vrf/regTable[2][6] , \vrf/regTable[2][7] ,
         \vrf/regTable[2][8] , \vrf/regTable[2][9] , \vrf/regTable[2][10] ,
         \vrf/regTable[2][11] , \vrf/regTable[2][12] , \vrf/regTable[2][13] ,
         \vrf/regTable[2][14] , \vrf/regTable[2][15] , \vrf/regTable[2][16] ,
         \vrf/regTable[2][17] , \vrf/regTable[2][18] , \vrf/regTable[2][19] ,
         \vrf/regTable[2][20] , \vrf/regTable[2][21] , \vrf/regTable[2][22] ,
         \vrf/regTable[2][23] , \vrf/regTable[2][24] , \vrf/regTable[2][25] ,
         \vrf/regTable[2][26] , \vrf/regTable[2][27] , \vrf/regTable[2][28] ,
         \vrf/regTable[2][29] , \vrf/regTable[2][30] , \vrf/regTable[2][31] ,
         \vrf/regTable[2][32] , \vrf/regTable[2][33] , \vrf/regTable[2][34] ,
         \vrf/regTable[2][35] , \vrf/regTable[2][36] , \vrf/regTable[2][37] ,
         \vrf/regTable[2][38] , \vrf/regTable[2][39] , \vrf/regTable[2][40] ,
         \vrf/regTable[2][41] , \vrf/regTable[2][42] , \vrf/regTable[2][43] ,
         \vrf/regTable[2][44] , \vrf/regTable[2][45] , \vrf/regTable[2][46] ,
         \vrf/regTable[2][47] , \vrf/regTable[2][48] , \vrf/regTable[2][49] ,
         \vrf/regTable[2][50] , \vrf/regTable[2][51] , \vrf/regTable[2][52] ,
         \vrf/regTable[2][53] , \vrf/regTable[2][54] , \vrf/regTable[2][55] ,
         \vrf/regTable[2][56] , \vrf/regTable[2][57] , \vrf/regTable[2][58] ,
         \vrf/regTable[2][59] , \vrf/regTable[2][60] , \vrf/regTable[2][61] ,
         \vrf/regTable[2][62] , \vrf/regTable[2][63] , \vrf/regTable[2][64] ,
         \vrf/regTable[2][65] , \vrf/regTable[2][66] , \vrf/regTable[2][67] ,
         \vrf/regTable[2][68] , \vrf/regTable[2][69] , \vrf/regTable[2][70] ,
         \vrf/regTable[2][71] , \vrf/regTable[2][72] , \vrf/regTable[2][73] ,
         \vrf/regTable[2][74] , \vrf/regTable[2][75] , \vrf/regTable[2][76] ,
         \vrf/regTable[2][77] , \vrf/regTable[2][78] , \vrf/regTable[2][79] ,
         \vrf/regTable[2][80] , \vrf/regTable[2][81] , \vrf/regTable[2][82] ,
         \vrf/regTable[2][83] , \vrf/regTable[2][84] , \vrf/regTable[2][85] ,
         \vrf/regTable[2][86] , \vrf/regTable[2][87] , \vrf/regTable[2][88] ,
         \vrf/regTable[2][89] , \vrf/regTable[2][90] , \vrf/regTable[2][91] ,
         \vrf/regTable[2][92] , \vrf/regTable[2][93] , \vrf/regTable[2][94] ,
         \vrf/regTable[2][95] , \vrf/regTable[2][96] , \vrf/regTable[2][97] ,
         \vrf/regTable[2][98] , \vrf/regTable[2][99] , \vrf/regTable[2][100] ,
         \vrf/regTable[2][101] , \vrf/regTable[2][102] ,
         \vrf/regTable[2][103] , \vrf/regTable[2][104] ,
         \vrf/regTable[2][105] , \vrf/regTable[2][106] ,
         \vrf/regTable[2][107] , \vrf/regTable[2][108] ,
         \vrf/regTable[2][109] , \vrf/regTable[2][110] ,
         \vrf/regTable[2][111] , \vrf/regTable[2][112] ,
         \vrf/regTable[2][113] , \vrf/regTable[2][114] ,
         \vrf/regTable[2][115] , \vrf/regTable[2][116] ,
         \vrf/regTable[2][117] , \vrf/regTable[2][118] ,
         \vrf/regTable[2][119] , \vrf/regTable[2][120] ,
         \vrf/regTable[2][121] , \vrf/regTable[2][122] ,
         \vrf/regTable[2][123] , \vrf/regTable[2][124] ,
         \vrf/regTable[2][125] , \vrf/regTable[2][126] ,
         \vrf/regTable[2][127] , \vrf/regTable[2][128] ,
         \vrf/regTable[2][129] , \vrf/regTable[2][130] ,
         \vrf/regTable[2][131] , \vrf/regTable[2][132] ,
         \vrf/regTable[2][133] , \vrf/regTable[2][134] ,
         \vrf/regTable[2][135] , \vrf/regTable[2][136] ,
         \vrf/regTable[2][137] , \vrf/regTable[2][138] ,
         \vrf/regTable[2][139] , \vrf/regTable[2][140] ,
         \vrf/regTable[2][141] , \vrf/regTable[2][142] ,
         \vrf/regTable[2][143] , \vrf/regTable[2][144] ,
         \vrf/regTable[2][145] , \vrf/regTable[2][146] ,
         \vrf/regTable[2][147] , \vrf/regTable[2][148] ,
         \vrf/regTable[2][149] , \vrf/regTable[2][150] ,
         \vrf/regTable[2][151] , \vrf/regTable[2][152] ,
         \vrf/regTable[2][153] , \vrf/regTable[2][154] ,
         \vrf/regTable[2][155] , \vrf/regTable[2][156] ,
         \vrf/regTable[2][157] , \vrf/regTable[2][158] ,
         \vrf/regTable[2][159] , \vrf/regTable[2][160] ,
         \vrf/regTable[2][161] , \vrf/regTable[2][162] ,
         \vrf/regTable[2][163] , \vrf/regTable[2][164] ,
         \vrf/regTable[2][165] , \vrf/regTable[2][166] ,
         \vrf/regTable[2][167] , \vrf/regTable[2][168] ,
         \vrf/regTable[2][169] , \vrf/regTable[2][170] ,
         \vrf/regTable[2][171] , \vrf/regTable[2][172] ,
         \vrf/regTable[2][173] , \vrf/regTable[2][174] ,
         \vrf/regTable[2][175] , \vrf/regTable[2][176] ,
         \vrf/regTable[2][177] , \vrf/regTable[2][178] ,
         \vrf/regTable[2][179] , \vrf/regTable[2][180] ,
         \vrf/regTable[2][181] , \vrf/regTable[2][182] ,
         \vrf/regTable[2][183] , \vrf/regTable[2][184] ,
         \vrf/regTable[2][185] , \vrf/regTable[2][186] ,
         \vrf/regTable[2][187] , \vrf/regTable[2][188] ,
         \vrf/regTable[2][189] , \vrf/regTable[2][190] ,
         \vrf/regTable[2][191] , \vrf/regTable[2][192] ,
         \vrf/regTable[2][193] , \vrf/regTable[2][194] ,
         \vrf/regTable[2][195] , \vrf/regTable[2][196] ,
         \vrf/regTable[2][197] , \vrf/regTable[2][198] ,
         \vrf/regTable[2][199] , \vrf/regTable[2][200] ,
         \vrf/regTable[2][201] , \vrf/regTable[2][202] ,
         \vrf/regTable[2][203] , \vrf/regTable[2][204] ,
         \vrf/regTable[2][205] , \vrf/regTable[2][206] ,
         \vrf/regTable[2][207] , \vrf/regTable[2][208] ,
         \vrf/regTable[2][209] , \vrf/regTable[2][210] ,
         \vrf/regTable[2][211] , \vrf/regTable[2][212] ,
         \vrf/regTable[2][213] , \vrf/regTable[2][214] ,
         \vrf/regTable[2][215] , \vrf/regTable[2][216] ,
         \vrf/regTable[2][217] , \vrf/regTable[2][218] ,
         \vrf/regTable[2][219] , \vrf/regTable[2][220] ,
         \vrf/regTable[2][221] , \vrf/regTable[2][222] ,
         \vrf/regTable[2][223] , \vrf/regTable[2][224] ,
         \vrf/regTable[2][225] , \vrf/regTable[2][226] ,
         \vrf/regTable[2][227] , \vrf/regTable[2][228] ,
         \vrf/regTable[2][229] , \vrf/regTable[2][230] ,
         \vrf/regTable[2][231] , \vrf/regTable[2][232] ,
         \vrf/regTable[2][233] , \vrf/regTable[2][234] ,
         \vrf/regTable[2][235] , \vrf/regTable[2][236] ,
         \vrf/regTable[2][237] , \vrf/regTable[2][238] ,
         \vrf/regTable[2][239] , \vrf/regTable[2][240] ,
         \vrf/regTable[2][241] , \vrf/regTable[2][242] ,
         \vrf/regTable[2][243] , \vrf/regTable[2][244] ,
         \vrf/regTable[2][245] , \vrf/regTable[2][246] ,
         \vrf/regTable[2][247] , \vrf/regTable[2][248] ,
         \vrf/regTable[2][249] , \vrf/regTable[2][250] ,
         \vrf/regTable[2][251] , \vrf/regTable[2][252] ,
         \vrf/regTable[2][253] , \vrf/regTable[2][254] ,
         \vrf/regTable[2][255] , \vrf/regTable[1][0] , \vrf/regTable[1][1] ,
         \vrf/regTable[1][2] , \vrf/regTable[1][3] , \vrf/regTable[1][4] ,
         \vrf/regTable[1][5] , \vrf/regTable[1][6] , \vrf/regTable[1][7] ,
         \vrf/regTable[1][8] , \vrf/regTable[1][9] , \vrf/regTable[1][10] ,
         \vrf/regTable[1][11] , \vrf/regTable[1][12] , \vrf/regTable[1][13] ,
         \vrf/regTable[1][14] , \vrf/regTable[1][15] , \vrf/regTable[1][16] ,
         \vrf/regTable[1][17] , \vrf/regTable[1][18] , \vrf/regTable[1][19] ,
         \vrf/regTable[1][20] , \vrf/regTable[1][21] , \vrf/regTable[1][22] ,
         \vrf/regTable[1][23] , \vrf/regTable[1][24] , \vrf/regTable[1][25] ,
         \vrf/regTable[1][26] , \vrf/regTable[1][27] , \vrf/regTable[1][28] ,
         \vrf/regTable[1][29] , \vrf/regTable[1][30] , \vrf/regTable[1][31] ,
         \vrf/regTable[1][32] , \vrf/regTable[1][33] , \vrf/regTable[1][34] ,
         \vrf/regTable[1][35] , \vrf/regTable[1][36] , \vrf/regTable[1][37] ,
         \vrf/regTable[1][38] , \vrf/regTable[1][39] , \vrf/regTable[1][40] ,
         \vrf/regTable[1][41] , \vrf/regTable[1][42] , \vrf/regTable[1][43] ,
         \vrf/regTable[1][44] , \vrf/regTable[1][45] , \vrf/regTable[1][46] ,
         \vrf/regTable[1][47] , \vrf/regTable[1][48] , \vrf/regTable[1][49] ,
         \vrf/regTable[1][50] , \vrf/regTable[1][51] , \vrf/regTable[1][52] ,
         \vrf/regTable[1][53] , \vrf/regTable[1][54] , \vrf/regTable[1][55] ,
         \vrf/regTable[1][56] , \vrf/regTable[1][57] , \vrf/regTable[1][58] ,
         \vrf/regTable[1][59] , \vrf/regTable[1][60] , \vrf/regTable[1][61] ,
         \vrf/regTable[1][62] , \vrf/regTable[1][63] , \vrf/regTable[1][64] ,
         \vrf/regTable[1][65] , \vrf/regTable[1][66] , \vrf/regTable[1][67] ,
         \vrf/regTable[1][68] , \vrf/regTable[1][69] , \vrf/regTable[1][70] ,
         \vrf/regTable[1][71] , \vrf/regTable[1][72] , \vrf/regTable[1][73] ,
         \vrf/regTable[1][74] , \vrf/regTable[1][75] , \vrf/regTable[1][76] ,
         \vrf/regTable[1][77] , \vrf/regTable[1][78] , \vrf/regTable[1][79] ,
         \vrf/regTable[1][80] , \vrf/regTable[1][81] , \vrf/regTable[1][82] ,
         \vrf/regTable[1][83] , \vrf/regTable[1][84] , \vrf/regTable[1][85] ,
         \vrf/regTable[1][86] , \vrf/regTable[1][87] , \vrf/regTable[1][88] ,
         \vrf/regTable[1][89] , \vrf/regTable[1][90] , \vrf/regTable[1][91] ,
         \vrf/regTable[1][92] , \vrf/regTable[1][93] , \vrf/regTable[1][94] ,
         \vrf/regTable[1][95] , \vrf/regTable[1][96] , \vrf/regTable[1][97] ,
         \vrf/regTable[1][98] , \vrf/regTable[1][99] , \vrf/regTable[1][100] ,
         \vrf/regTable[1][101] , \vrf/regTable[1][102] ,
         \vrf/regTable[1][103] , \vrf/regTable[1][104] ,
         \vrf/regTable[1][105] , \vrf/regTable[1][106] ,
         \vrf/regTable[1][107] , \vrf/regTable[1][108] ,
         \vrf/regTable[1][109] , \vrf/regTable[1][110] ,
         \vrf/regTable[1][111] , \vrf/regTable[1][112] ,
         \vrf/regTable[1][113] , \vrf/regTable[1][114] ,
         \vrf/regTable[1][115] , \vrf/regTable[1][116] ,
         \vrf/regTable[1][117] , \vrf/regTable[1][118] ,
         \vrf/regTable[1][119] , \vrf/regTable[1][120] ,
         \vrf/regTable[1][121] , \vrf/regTable[1][122] ,
         \vrf/regTable[1][123] , \vrf/regTable[1][124] ,
         \vrf/regTable[1][125] , \vrf/regTable[1][126] ,
         \vrf/regTable[1][127] , \vrf/regTable[1][128] ,
         \vrf/regTable[1][129] , \vrf/regTable[1][130] ,
         \vrf/regTable[1][131] , \vrf/regTable[1][132] ,
         \vrf/regTable[1][133] , \vrf/regTable[1][134] ,
         \vrf/regTable[1][135] , \vrf/regTable[1][136] ,
         \vrf/regTable[1][137] , \vrf/regTable[1][138] ,
         \vrf/regTable[1][139] , \vrf/regTable[1][140] ,
         \vrf/regTable[1][141] , \vrf/regTable[1][142] ,
         \vrf/regTable[1][143] , \vrf/regTable[1][144] ,
         \vrf/regTable[1][145] , \vrf/regTable[1][146] ,
         \vrf/regTable[1][147] , \vrf/regTable[1][148] ,
         \vrf/regTable[1][149] , \vrf/regTable[1][150] ,
         \vrf/regTable[1][151] , \vrf/regTable[1][152] ,
         \vrf/regTable[1][153] , \vrf/regTable[1][154] ,
         \vrf/regTable[1][155] , \vrf/regTable[1][156] ,
         \vrf/regTable[1][157] , \vrf/regTable[1][158] ,
         \vrf/regTable[1][159] , \vrf/regTable[1][160] ,
         \vrf/regTable[1][161] , \vrf/regTable[1][162] ,
         \vrf/regTable[1][163] , \vrf/regTable[1][164] ,
         \vrf/regTable[1][165] , \vrf/regTable[1][166] ,
         \vrf/regTable[1][167] , \vrf/regTable[1][168] ,
         \vrf/regTable[1][169] , \vrf/regTable[1][170] ,
         \vrf/regTable[1][171] , \vrf/regTable[1][172] ,
         \vrf/regTable[1][173] , \vrf/regTable[1][174] ,
         \vrf/regTable[1][175] , \vrf/regTable[1][176] ,
         \vrf/regTable[1][177] , \vrf/regTable[1][178] ,
         \vrf/regTable[1][179] , \vrf/regTable[1][180] ,
         \vrf/regTable[1][181] , \vrf/regTable[1][182] ,
         \vrf/regTable[1][183] , \vrf/regTable[1][184] ,
         \vrf/regTable[1][185] , \vrf/regTable[1][186] ,
         \vrf/regTable[1][187] , \vrf/regTable[1][188] ,
         \vrf/regTable[1][189] , \vrf/regTable[1][190] ,
         \vrf/regTable[1][191] , \vrf/regTable[1][192] ,
         \vrf/regTable[1][193] , \vrf/regTable[1][194] ,
         \vrf/regTable[1][195] , \vrf/regTable[1][196] ,
         \vrf/regTable[1][197] , \vrf/regTable[1][198] ,
         \vrf/regTable[1][199] , \vrf/regTable[1][200] ,
         \vrf/regTable[1][201] , \vrf/regTable[1][202] ,
         \vrf/regTable[1][203] , \vrf/regTable[1][204] ,
         \vrf/regTable[1][205] , \vrf/regTable[1][206] ,
         \vrf/regTable[1][207] , \vrf/regTable[1][208] ,
         \vrf/regTable[1][209] , \vrf/regTable[1][210] ,
         \vrf/regTable[1][211] , \vrf/regTable[1][212] ,
         \vrf/regTable[1][213] , \vrf/regTable[1][214] ,
         \vrf/regTable[1][215] , \vrf/regTable[1][216] ,
         \vrf/regTable[1][217] , \vrf/regTable[1][218] ,
         \vrf/regTable[1][219] , \vrf/regTable[1][220] ,
         \vrf/regTable[1][221] , \vrf/regTable[1][222] ,
         \vrf/regTable[1][223] , \vrf/regTable[1][224] ,
         \vrf/regTable[1][225] , \vrf/regTable[1][226] ,
         \vrf/regTable[1][227] , \vrf/regTable[1][228] ,
         \vrf/regTable[1][229] , \vrf/regTable[1][230] ,
         \vrf/regTable[1][231] , \vrf/regTable[1][232] ,
         \vrf/regTable[1][233] , \vrf/regTable[1][234] ,
         \vrf/regTable[1][235] , \vrf/regTable[1][236] ,
         \vrf/regTable[1][237] , \vrf/regTable[1][238] ,
         \vrf/regTable[1][239] , \vrf/regTable[1][240] ,
         \vrf/regTable[1][241] , \vrf/regTable[1][242] ,
         \vrf/regTable[1][243] , \vrf/regTable[1][244] ,
         \vrf/regTable[1][245] , \vrf/regTable[1][246] ,
         \vrf/regTable[1][247] , \vrf/regTable[1][248] ,
         \vrf/regTable[1][249] , \vrf/regTable[1][250] ,
         \vrf/regTable[1][251] , \vrf/regTable[1][252] ,
         \vrf/regTable[1][253] , \vrf/regTable[1][254] ,
         \vrf/regTable[1][255] , \vrf/regTable[0][0] , \vrf/regTable[0][1] ,
         \vrf/regTable[0][2] , \vrf/regTable[0][3] , \vrf/regTable[0][4] ,
         \vrf/regTable[0][5] , \vrf/regTable[0][6] , \vrf/regTable[0][7] ,
         \vrf/regTable[0][8] , \vrf/regTable[0][9] , \vrf/regTable[0][10] ,
         \vrf/regTable[0][11] , \vrf/regTable[0][12] , \vrf/regTable[0][13] ,
         \vrf/regTable[0][14] , \vrf/regTable[0][15] , \vrf/regTable[0][16] ,
         \vrf/regTable[0][17] , \vrf/regTable[0][18] , \vrf/regTable[0][19] ,
         \vrf/regTable[0][20] , \vrf/regTable[0][21] , \vrf/regTable[0][22] ,
         \vrf/regTable[0][23] , \vrf/regTable[0][24] , \vrf/regTable[0][25] ,
         \vrf/regTable[0][26] , \vrf/regTable[0][27] , \vrf/regTable[0][28] ,
         \vrf/regTable[0][29] , \vrf/regTable[0][30] , \vrf/regTable[0][31] ,
         \vrf/regTable[0][32] , \vrf/regTable[0][33] , \vrf/regTable[0][34] ,
         \vrf/regTable[0][35] , \vrf/regTable[0][36] , \vrf/regTable[0][37] ,
         \vrf/regTable[0][38] , \vrf/regTable[0][39] , \vrf/regTable[0][40] ,
         \vrf/regTable[0][41] , \vrf/regTable[0][42] , \vrf/regTable[0][43] ,
         \vrf/regTable[0][44] , \vrf/regTable[0][45] , \vrf/regTable[0][46] ,
         \vrf/regTable[0][47] , \vrf/regTable[0][48] , \vrf/regTable[0][49] ,
         \vrf/regTable[0][50] , \vrf/regTable[0][51] , \vrf/regTable[0][52] ,
         \vrf/regTable[0][53] , \vrf/regTable[0][54] , \vrf/regTable[0][55] ,
         \vrf/regTable[0][56] , \vrf/regTable[0][57] , \vrf/regTable[0][58] ,
         \vrf/regTable[0][59] , \vrf/regTable[0][60] , \vrf/regTable[0][61] ,
         \vrf/regTable[0][62] , \vrf/regTable[0][63] , \vrf/regTable[0][64] ,
         \vrf/regTable[0][65] , \vrf/regTable[0][66] , \vrf/regTable[0][67] ,
         \vrf/regTable[0][68] , \vrf/regTable[0][69] , \vrf/regTable[0][70] ,
         \vrf/regTable[0][71] , \vrf/regTable[0][72] , \vrf/regTable[0][73] ,
         \vrf/regTable[0][74] , \vrf/regTable[0][75] , \vrf/regTable[0][76] ,
         \vrf/regTable[0][77] , \vrf/regTable[0][78] , \vrf/regTable[0][79] ,
         \vrf/regTable[0][80] , \vrf/regTable[0][81] , \vrf/regTable[0][82] ,
         \vrf/regTable[0][83] , \vrf/regTable[0][84] , \vrf/regTable[0][85] ,
         \vrf/regTable[0][86] , \vrf/regTable[0][87] , \vrf/regTable[0][88] ,
         \vrf/regTable[0][89] , \vrf/regTable[0][90] , \vrf/regTable[0][91] ,
         \vrf/regTable[0][92] , \vrf/regTable[0][93] , \vrf/regTable[0][94] ,
         \vrf/regTable[0][95] , \vrf/regTable[0][96] , \vrf/regTable[0][97] ,
         \vrf/regTable[0][98] , \vrf/regTable[0][99] , \vrf/regTable[0][100] ,
         \vrf/regTable[0][101] , \vrf/regTable[0][102] ,
         \vrf/regTable[0][103] , \vrf/regTable[0][104] ,
         \vrf/regTable[0][105] , \vrf/regTable[0][106] ,
         \vrf/regTable[0][107] , \vrf/regTable[0][108] ,
         \vrf/regTable[0][109] , \vrf/regTable[0][110] ,
         \vrf/regTable[0][111] , \vrf/regTable[0][112] ,
         \vrf/regTable[0][113] , \vrf/regTable[0][114] ,
         \vrf/regTable[0][115] , \vrf/regTable[0][116] ,
         \vrf/regTable[0][117] , \vrf/regTable[0][118] ,
         \vrf/regTable[0][119] , \vrf/regTable[0][120] ,
         \vrf/regTable[0][121] , \vrf/regTable[0][122] ,
         \vrf/regTable[0][123] , \vrf/regTable[0][124] ,
         \vrf/regTable[0][125] , \vrf/regTable[0][126] ,
         \vrf/regTable[0][127] , \vrf/regTable[0][128] ,
         \vrf/regTable[0][129] , \vrf/regTable[0][130] ,
         \vrf/regTable[0][131] , \vrf/regTable[0][132] ,
         \vrf/regTable[0][133] , \vrf/regTable[0][134] ,
         \vrf/regTable[0][135] , \vrf/regTable[0][136] ,
         \vrf/regTable[0][137] , \vrf/regTable[0][138] ,
         \vrf/regTable[0][139] , \vrf/regTable[0][140] ,
         \vrf/regTable[0][141] , \vrf/regTable[0][142] ,
         \vrf/regTable[0][143] , \vrf/regTable[0][144] ,
         \vrf/regTable[0][145] , \vrf/regTable[0][146] ,
         \vrf/regTable[0][147] , \vrf/regTable[0][148] ,
         \vrf/regTable[0][149] , \vrf/regTable[0][150] ,
         \vrf/regTable[0][151] , \vrf/regTable[0][152] ,
         \vrf/regTable[0][153] , \vrf/regTable[0][154] ,
         \vrf/regTable[0][155] , \vrf/regTable[0][156] ,
         \vrf/regTable[0][157] , \vrf/regTable[0][158] ,
         \vrf/regTable[0][159] , \vrf/regTable[0][160] ,
         \vrf/regTable[0][161] , \vrf/regTable[0][162] ,
         \vrf/regTable[0][163] , \vrf/regTable[0][164] ,
         \vrf/regTable[0][165] , \vrf/regTable[0][166] ,
         \vrf/regTable[0][167] , \vrf/regTable[0][168] ,
         \vrf/regTable[0][169] , \vrf/regTable[0][170] ,
         \vrf/regTable[0][171] , \vrf/regTable[0][172] ,
         \vrf/regTable[0][173] , \vrf/regTable[0][174] ,
         \vrf/regTable[0][175] , \vrf/regTable[0][176] ,
         \vrf/regTable[0][177] , \vrf/regTable[0][178] ,
         \vrf/regTable[0][179] , \vrf/regTable[0][180] ,
         \vrf/regTable[0][181] , \vrf/regTable[0][182] ,
         \vrf/regTable[0][183] , \vrf/regTable[0][184] ,
         \vrf/regTable[0][185] , \vrf/regTable[0][186] ,
         \vrf/regTable[0][187] , \vrf/regTable[0][188] ,
         \vrf/regTable[0][189] , \vrf/regTable[0][190] ,
         \vrf/regTable[0][191] , \vrf/regTable[0][192] ,
         \vrf/regTable[0][193] , \vrf/regTable[0][194] ,
         \vrf/regTable[0][195] , \vrf/regTable[0][196] ,
         \vrf/regTable[0][197] , \vrf/regTable[0][198] ,
         \vrf/regTable[0][199] , \vrf/regTable[0][200] ,
         \vrf/regTable[0][201] , \vrf/regTable[0][202] ,
         \vrf/regTable[0][203] , \vrf/regTable[0][204] ,
         \vrf/regTable[0][205] , \vrf/regTable[0][206] ,
         \vrf/regTable[0][207] , \vrf/regTable[0][208] ,
         \vrf/regTable[0][209] , \vrf/regTable[0][210] ,
         \vrf/regTable[0][211] , \vrf/regTable[0][212] ,
         \vrf/regTable[0][213] , \vrf/regTable[0][214] ,
         \vrf/regTable[0][215] , \vrf/regTable[0][216] ,
         \vrf/regTable[0][217] , \vrf/regTable[0][218] ,
         \vrf/regTable[0][219] , \vrf/regTable[0][220] ,
         \vrf/regTable[0][221] , \vrf/regTable[0][222] ,
         \vrf/regTable[0][223] , \vrf/regTable[0][224] ,
         \vrf/regTable[0][225] , \vrf/regTable[0][226] ,
         \vrf/regTable[0][227] , \vrf/regTable[0][228] ,
         \vrf/regTable[0][229] , \vrf/regTable[0][230] ,
         \vrf/regTable[0][231] , \vrf/regTable[0][232] ,
         \vrf/regTable[0][233] , \vrf/regTable[0][234] ,
         \vrf/regTable[0][235] , \vrf/regTable[0][236] ,
         \vrf/regTable[0][237] , \vrf/regTable[0][238] ,
         \vrf/regTable[0][239] , \vrf/regTable[0][240] ,
         \vrf/regTable[0][241] , \vrf/regTable[0][242] ,
         \vrf/regTable[0][243] , \vrf/regTable[0][244] ,
         \vrf/regTable[0][245] , \vrf/regTable[0][246] ,
         \vrf/regTable[0][247] , \vrf/regTable[0][248] ,
         \vrf/regTable[0][249] , \vrf/regTable[0][250] ,
         \vrf/regTable[0][251] , \vrf/regTable[0][252] ,
         \vrf/regTable[0][253] , \vrf/regTable[0][254] ,
         \vrf/regTable[0][255] , \vrf/N14 , \vrf/N13 , \vrf/N12 , \vrf/N11 ,
         \vrf/N10 , \vrf/N9 , \srf/N59 , \srf/N58 , \srf/N57 , \srf/N56 ,
         \srf/N55 , \srf/N54 , \srf/N53 , \srf/N52 , \srf/N51 , \srf/N50 ,
         \srf/N49 , \srf/N48 , \srf/N47 , \srf/N46 , \srf/N45 , \srf/N44 ,
         \srf/N43 , \srf/N42 , \srf/N41 , \srf/N40 , \srf/N39 , \srf/N38 ,
         \srf/N37 , \srf/N36 , \srf/N35 , \srf/N34 , \srf/N33 , \srf/N32 ,
         \srf/N31 , \srf/N30 , \srf/N29 , \srf/N28 , \srf/N27 , \srf/N26 ,
         \srf/N25 , \srf/N24 , \srf/N23 , \srf/N22 , \srf/N21 , \srf/N20 ,
         \srf/regTable[7][0] , \srf/regTable[7][1] , \srf/regTable[7][2] ,
         \srf/regTable[7][3] , \srf/regTable[7][4] , \srf/regTable[7][5] ,
         \srf/regTable[7][6] , \srf/regTable[7][7] , \srf/regTable[7][8] ,
         \srf/regTable[7][9] , \srf/regTable[7][10] , \srf/regTable[7][11] ,
         \srf/regTable[7][12] , \srf/regTable[7][13] , \srf/regTable[7][14] ,
         \srf/regTable[7][15] , \srf/regTable[6][0] , \srf/regTable[6][1] ,
         \srf/regTable[6][2] , \srf/regTable[6][3] , \srf/regTable[6][4] ,
         \srf/regTable[6][5] , \srf/regTable[6][6] , \srf/regTable[6][7] ,
         \srf/regTable[6][8] , \srf/regTable[6][9] , \srf/regTable[6][10] ,
         \srf/regTable[6][11] , \srf/regTable[6][12] , \srf/regTable[6][13] ,
         \srf/regTable[6][14] , \srf/regTable[6][15] , \srf/regTable[5][0] ,
         \srf/regTable[5][1] , \srf/regTable[5][2] , \srf/regTable[5][3] ,
         \srf/regTable[5][4] , \srf/regTable[5][5] , \srf/regTable[5][6] ,
         \srf/regTable[5][7] , \srf/regTable[5][8] , \srf/regTable[5][9] ,
         \srf/regTable[5][10] , \srf/regTable[5][11] , \srf/regTable[5][12] ,
         \srf/regTable[5][13] , \srf/regTable[5][14] , \srf/regTable[5][15] ,
         \srf/regTable[4][0] , \srf/regTable[4][1] , \srf/regTable[4][2] ,
         \srf/regTable[4][3] , \srf/regTable[4][4] , \srf/regTable[4][5] ,
         \srf/regTable[4][6] , \srf/regTable[4][7] , \srf/regTable[4][8] ,
         \srf/regTable[4][9] , \srf/regTable[4][10] , \srf/regTable[4][11] ,
         \srf/regTable[4][12] , \srf/regTable[4][13] , \srf/regTable[4][14] ,
         \srf/regTable[4][15] , \srf/regTable[3][0] , \srf/regTable[3][1] ,
         \srf/regTable[3][2] , \srf/regTable[3][3] , \srf/regTable[3][4] ,
         \srf/regTable[3][5] , \srf/regTable[3][6] , \srf/regTable[3][7] ,
         \srf/regTable[3][8] , \srf/regTable[3][9] , \srf/regTable[3][10] ,
         \srf/regTable[3][11] , \srf/regTable[3][12] , \srf/regTable[3][13] ,
         \srf/regTable[3][14] , \srf/regTable[3][15] , \srf/regTable[2][0] ,
         \srf/regTable[2][1] , \srf/regTable[2][2] , \srf/regTable[2][3] ,
         \srf/regTable[2][4] , \srf/regTable[2][5] , \srf/regTable[2][6] ,
         \srf/regTable[2][7] , \srf/regTable[2][8] , \srf/regTable[2][9] ,
         \srf/regTable[2][10] , \srf/regTable[2][11] , \srf/regTable[2][12] ,
         \srf/regTable[2][13] , \srf/regTable[2][14] , \srf/regTable[2][15] ,
         \srf/regTable[1][0] , \srf/regTable[1][1] , \srf/regTable[1][2] ,
         \srf/regTable[1][3] , \srf/regTable[1][4] , \srf/regTable[1][5] ,
         \srf/regTable[1][6] , \srf/regTable[1][7] , \srf/regTable[1][8] ,
         \srf/regTable[1][9] , \srf/regTable[1][10] , \srf/regTable[1][11] ,
         \srf/regTable[1][12] , \srf/regTable[1][13] , \srf/regTable[1][14] ,
         \srf/regTable[1][15] , \srf/regTable[0][0] , \srf/regTable[0][1] ,
         \srf/regTable[0][2] , \srf/regTable[0][3] , \srf/regTable[0][4] ,
         \srf/regTable[0][5] , \srf/regTable[0][6] , \srf/regTable[0][7] ,
         \srf/regTable[0][8] , \srf/regTable[0][9] , \srf/regTable[0][10] ,
         \srf/regTable[0][11] , \srf/regTable[0][12] , \srf/regTable[0][13] ,
         \srf/regTable[0][14] , \srf/regTable[0][15] , \srf/N17 , \srf/N15 ,
         \alu/N1019 , \alu/N1018 , \alu/N1016 , \alu/N1015 , \alu/N1014 ,
         \alu/N1011 , \alu/N1003 , \alu/N990 , \alu/N989 , \alu/N988 ,
         \alu/N986 , \alu/N984 , \alu/N983 , \alu/N832 , \alu/N808 ,
         \alu/N684 , \alu/N683 , \alu/N665 , \alu/N661 , \alu/N659 ,
         \alu/N657 , \alu/N655 , \alu/N653 , \alu/N634 , \alu/N339 ,
         \alu/N338 , \alu/N337 , \alu/N336 , \alu/N335 , \alu/N334 ,
         \alu/N333 , \alu/N332 , \alu/N331 , \alu/N330 , \alu/N329 ,
         \alu/N328 , \alu/N327 , \alu/N326 , \alu/N325 , \alu/N324 ,
         \alu/N323 , \alu/N322 , \alu/N321 , \alu/N320 , \alu/N319 ,
         \alu/N318 , \alu/N317 , \alu/N316 , \alu/N315 , \alu/N314 ,
         \alu/N313 , \alu/N88 , \alu/N87 , n1, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n132, n134, n136, n137, n138, n153, n156, n3020, \mult_x_153/n181 ,
         \mult_x_153/n180 , \mult_x_153/n179 , \mult_x_153/n178 ,
         \mult_x_153/n177 , \mult_x_153/n176 , \mult_x_153/n170 ,
         \mult_x_153/n169 , \mult_x_153/n168 , \mult_x_153/n166 ,
         \mult_x_153/n165 , \mult_x_153/n164 , \mult_x_153/n163 ,
         \mult_x_153/n162 , \mult_x_153/n159 , \mult_x_153/n158 ,
         \mult_x_153/n155 , \mult_x_153/n154 , \mult_x_153/n153 ,
         \mult_x_153/n152 , \mult_x_153/n151 , \mult_x_153/n150 ,
         \mult_x_153/n149 , \mult_x_153/n148 , \mult_x_153/n144 ,
         \mult_x_153/n143 , \mult_x_153/n142 , \mult_x_153/n141 ,
         \mult_x_153/n140 , \mult_x_153/n137 , \mult_x_153/n136 ,
         \mult_x_153/n133 , \mult_x_153/n132 , \mult_x_153/n131 ,
         \mult_x_153/n130 , \mult_x_153/n129 , \mult_x_153/n127 ,
         \mult_x_153/n126 , \mult_x_153/n125 , \mult_x_153/n122 ,
         \mult_x_153/n121 , \mult_x_153/n120 , \mult_x_153/n119 ,
         \mult_x_153/n117 , \mult_x_153/n105 , \mult_x_153/n102 ,
         \mult_x_153/n101 , \mult_x_153/n100 , \mult_x_153/n99 ,
         \mult_x_153/n98 , \mult_x_153/n97 , \mult_x_153/n96 ,
         \mult_x_153/n95 , \mult_x_153/n94 , \mult_x_153/n93 ,
         \mult_x_153/n92 , \mult_x_153/n91 , \mult_x_153/n90 ,
         \mult_x_153/n89 , \mult_x_153/n88 , \mult_x_153/n87 ,
         \mult_x_153/n86 , \mult_x_153/n85 , \mult_x_153/n84 ,
         \mult_x_153/n83 , \mult_x_153/n82 , \mult_x_153/n81 ,
         \mult_x_153/n80 , \mult_x_153/n79 , \mult_x_153/n78 ,
         \mult_x_153/n77 , \mult_x_153/n76 , \mult_x_153/n75 ,
         \mult_x_153/n74 , \mult_x_153/n73 , \mult_x_153/n72 ,
         \mult_x_153/n71 , \mult_x_153/n70 , \mult_x_153/n69 ,
         \mult_x_153/n68 , \mult_x_153/n67 , \mult_x_153/n66 ,
         \mult_x_153/n65 , \mult_x_153/n64 , \mult_x_153/n61 ,
         \mult_x_153/n60 , \mult_x_153/n59 , \mult_x_153/n58 ,
         \mult_x_153/n57 , \mult_x_153/n56 , \mult_x_153/n55 ,
         \mult_x_153/n54 , \mult_x_153/n53 , \mult_x_153/n52 ,
         \mult_x_153/n51 , \mult_x_153/n50 , \mult_x_153/n47 ,
         \mult_x_153/n46 , \mult_x_153/n45 , \mult_x_153/n44 ,
         \mult_x_153/n43 , \mult_x_153/n42 , \mult_x_153/n41 ,
         \mult_x_153/n40 , \mult_x_153/n39 , \mult_x_153/n38 ,
         \mult_x_153/n37 , \mult_x_153/n35 , \mult_x_153/n34 ,
         \mult_x_153/n33 , \mult_x_153/n32 , \mult_x_153/n31 ,
         \mult_x_153/n30 , \C1/Z_0 , \C2/Z_25 , \C2/Z_24 , \C2/Z_23 ,
         \C2/Z_22 , \C2/Z_21 , \C2/Z_20 , \C2/Z_19 , \C2/Z_18 , \C2/Z_17 ,
         \C2/Z_16 , \C3/Z_25 , \C3/Z_24 , \C3/Z_23 , \C3/Z_22 , \C3/Z_21 ,
         \C3/Z_19 , \C3/Z_18 , \C3/Z_17 , \C3/Z_16 , \C3/Z_14 , \C3/Z_13 ,
         \C3/Z_12 , \C3/Z_11 , \C3/Z_10 , \C3/Z_9 , \C3/Z_8 , \C3/Z_7 ,
         \C3/Z_6 , \C3/Z_5 , \C3/Z_4 , \C3/Z_3 , \C3/Z_2 , \C3/Z_1 , \C3/Z_0 ,
         \DP_OP_487J11_125_9213/n56 , \DP_OP_487J11_125_9213/n55 ,
         \DP_OP_487J11_125_9213/n54 , \DP_OP_487J11_125_9213/n53 ,
         \DP_OP_487J11_125_9213/n52 , \DP_OP_487J11_125_9213/n51 ,
         \DP_OP_487J11_125_9213/n50 , \DP_OP_487J11_125_9213/n49 ,
         \DP_OP_487J11_125_9213/n48 , \DP_OP_487J11_125_9213/n47 ,
         \DP_OP_487J11_125_9213/n46 , \DP_OP_487J11_125_9213/n45 ,
         \DP_OP_487J11_125_9213/n44 , \DP_OP_487J11_125_9213/n43 ,
         \DP_OP_487J11_125_9213/n42 , \DP_OP_487J11_125_9213/n40 ,
         \DP_OP_487J11_125_9213/n39 , \DP_OP_487J11_125_9213/n38 ,
         \DP_OP_487J11_125_9213/n37 , \DP_OP_487J11_125_9213/n36 ,
         \DP_OP_487J11_125_9213/n35 , \DP_OP_487J11_125_9213/n34 ,
         \DP_OP_487J11_125_9213/n33 , \DP_OP_487J11_125_9213/n32 ,
         \DP_OP_487J11_125_9213/n31 , \DP_OP_487J11_125_9213/n26 ,
         \DP_OP_487J11_125_9213/n25 , \DP_OP_487J11_125_9213/n24 ,
         \DP_OP_487J11_125_9213/n23 , \DP_OP_487J11_125_9213/n22 ,
         \DP_OP_487J11_125_9213/n21 , \DP_OP_487J11_125_9213/n20 ,
         \DP_OP_487J11_125_9213/n19 , \DP_OP_487J11_125_9213/n18 ,
         \DP_OP_487J11_125_9213/n17 , \DP_OP_487J11_125_9213/n16 ,
         \DP_OP_487J11_125_9213/n15 , \DP_OP_487J11_125_9213/n14 ,
         \DP_OP_487J11_125_9213/n13 , \DP_OP_487J11_125_9213/n11 ,
         \DP_OP_487J11_125_9213/n10 , \DP_OP_487J11_125_9213/n9 ,
         \DP_OP_487J11_125_9213/n8 , \DP_OP_487J11_125_9213/n7 ,
         \DP_OP_487J11_125_9213/n6 , \DP_OP_487J11_125_9213/n5 ,
         \DP_OP_487J11_125_9213/n4 , \DP_OP_487J11_125_9213/n3 ,
         \DP_OP_487J11_125_9213/n2 , \DP_OP_487J11_125_9213/n1 ,
         \DP_OP_493J11_130_7648/n56 , \DP_OP_493J11_130_7648/n55 ,
         \DP_OP_493J11_130_7648/n54 , \DP_OP_493J11_130_7648/n53 ,
         \DP_OP_493J11_130_7648/n52 , \DP_OP_493J11_130_7648/n51 ,
         \DP_OP_493J11_130_7648/n50 , \DP_OP_493J11_130_7648/n49 ,
         \DP_OP_493J11_130_7648/n48 , \DP_OP_493J11_130_7648/n47 ,
         \DP_OP_493J11_130_7648/n46 , \DP_OP_493J11_130_7648/n45 ,
         \DP_OP_493J11_130_7648/n44 , \DP_OP_493J11_130_7648/n43 ,
         \DP_OP_493J11_130_7648/n42 , \DP_OP_493J11_130_7648/n41 ,
         \DP_OP_493J11_130_7648/n40 , \DP_OP_493J11_130_7648/n39 ,
         \DP_OP_493J11_130_7648/n38 , \DP_OP_493J11_130_7648/n37 ,
         \DP_OP_493J11_130_7648/n36 , \DP_OP_493J11_130_7648/n35 ,
         \DP_OP_493J11_130_7648/n34 , \DP_OP_493J11_130_7648/n33 ,
         \DP_OP_493J11_130_7648/n32 , \DP_OP_493J11_130_7648/n31 ,
         \DP_OP_493J11_130_7648/n26 , \DP_OP_493J11_130_7648/n25 ,
         \DP_OP_493J11_130_7648/n24 , \DP_OP_493J11_130_7648/n23 ,
         \DP_OP_493J11_130_7648/n22 , \DP_OP_493J11_130_7648/n21 ,
         \DP_OP_493J11_130_7648/n20 , \DP_OP_493J11_130_7648/n19 ,
         \DP_OP_493J11_130_7648/n18 , \DP_OP_493J11_130_7648/n17 ,
         \DP_OP_493J11_130_7648/n16 , \DP_OP_493J11_130_7648/n15 ,
         \DP_OP_493J11_130_7648/n14 , \DP_OP_493J11_130_7648/n13 ,
         \DP_OP_493J11_130_7648/n12 , \DP_OP_493J11_130_7648/n11 ,
         \DP_OP_493J11_130_7648/n10 , \DP_OP_493J11_130_7648/n9 ,
         \DP_OP_493J11_130_7648/n8 , \DP_OP_493J11_130_7648/n7 ,
         \DP_OP_493J11_130_7648/n6 , \DP_OP_493J11_130_7648/n5 ,
         \DP_OP_493J11_130_7648/n4 , \DP_OP_493J11_130_7648/n3 ,
         \DP_OP_493J11_130_7648/n2 , \DP_OP_493J11_130_7648/n1 ,
         \intadd_33/A[9] , \intadd_33/B[9] , \intadd_33/B[8] , \intadd_33/CI ,
         \intadd_33/SUM[9] , \intadd_33/SUM[8] , \intadd_33/SUM[7] ,
         \intadd_33/SUM[6] , \intadd_33/SUM[5] , \intadd_33/SUM[4] ,
         \intadd_33/SUM[3] , \intadd_33/SUM[2] , \intadd_33/SUM[1] ,
         \intadd_33/SUM[0] , \intadd_33/n10 , \intadd_33/n9 , \intadd_33/n8 ,
         \intadd_33/n7 , \intadd_33/n6 , \intadd_33/n5 , \intadd_33/n4 ,
         \intadd_33/n3 , \intadd_33/n2 , \intadd_33/n1 , \intadd_34/A[3] ,
         \intadd_34/A[2] , \intadd_34/A[1] , \intadd_34/A[0] , \intadd_34/CI ,
         \intadd_34/SUM[3] , \intadd_34/SUM[2] , \intadd_34/SUM[1] ,
         \intadd_34/SUM[0] , \intadd_34/CO , \intadd_34/n4 , \intadd_34/n3 ,
         \intadd_34/n2 , \intadd_34/n1 , \intadd_35/A[2] , \intadd_35/A[1] ,
         \intadd_35/A[0] , \intadd_35/B[2] , \intadd_35/B[1] ,
         \intadd_35/B[0] , \intadd_35/CI , \intadd_35/SUM[2] ,
         \intadd_35/SUM[1] , \intadd_35/SUM[0] , \intadd_35/n3 ,
         \intadd_35/n2 , \intadd_35/n1 , \intadd_36/B[2] , \intadd_36/B[1] ,
         \intadd_36/B[0] , \intadd_36/CI , \intadd_36/SUM[2] ,
         \intadd_36/SUM[1] , \intadd_36/SUM[0] , \intadd_36/n3 ,
         \intadd_36/n2 , \intadd_36/n1 , n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4614,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336;
  wire   [255:0] vectorData1;
  wire   [255:0] vectorData2;
  wire   [15:0] scalarData1;
  wire   [15:0] scalarData2;
  wire   [255:0] op1;
  wire   [255:0] op2;
  wire   [3:0] func;
  wire   [255:0] result;
  wire   [15:0] instrIn;
  wire   [3:0] code;
  wire   [3:0] state;
  wire   [4:0] cycles;
  wire   [255:0] vectorToLoad;
  wire   [15:0] scalarToLoad;
  wire   [15:0] nextInstrAddr;

  LNQD1BWP \instrIn_reg[15]  ( .D(DataIn[15]), .EN(n3020), .Q(code[3]) );
  LNQD1BWP \instrIn_reg[14]  ( .D(DataIn[14]), .EN(n3020), .Q(code[2]) );
  LNQD1BWP \instrIn_reg[13]  ( .D(DataIn[13]), .EN(n3020), .Q(code[1]) );
  LHQD1BWP \func_reg[0]  ( .E(n4616), .D(code[0]), .Q(func[0]) );
  LHQD1BWP \func_reg[2]  ( .E(n4616), .D(code[2]), .Q(func[2]) );
  LHQD1BWP \func_reg[3]  ( .E(n4616), .D(code[3]), .Q(func[3]) );
  LHQD1BWP \scalarToLoad_reg[9]  ( .E(n4695), .D(N1819), .Q(scalarToLoad[9])
         );
  LHQD1BWP \scalarToLoad_reg[8]  ( .E(n4695), .D(N1818), .Q(scalarToLoad[8])
         );
  LHQD1BWP \scalarToLoad_reg[7]  ( .E(n4695), .D(N1817), .Q(scalarToLoad[7])
         );
  LHQD1BWP \scalarToLoad_reg[6]  ( .E(n4695), .D(N1816), .Q(scalarToLoad[6])
         );
  LHQD1BWP \scalarToLoad_reg[5]  ( .E(n4695), .D(N1815), .Q(scalarToLoad[5])
         );
  LHQD1BWP \scalarToLoad_reg[4]  ( .E(n4695), .D(N1814), .Q(scalarToLoad[4])
         );
  LHQD1BWP \scalarToLoad_reg[3]  ( .E(n4695), .D(N1813), .Q(scalarToLoad[3])
         );
  LHQD1BWP \scalarToLoad_reg[2]  ( .E(n4695), .D(N1812), .Q(scalarToLoad[2])
         );
  LHQD1BWP \scalarToLoad_reg[1]  ( .E(n4695), .D(N1811), .Q(scalarToLoad[1])
         );
  LHQD1BWP \scalarToLoad_reg[0]  ( .E(n4695), .D(N1810), .Q(scalarToLoad[0])
         );
  LHQD1BWP \scalarToLoad_reg[15]  ( .E(n4695), .D(N1825), .Q(scalarToLoad[15])
         );
  LHQD1BWP \nextInstrAddr_reg[9]  ( .E(N4162), .D(N4163), .Q(nextInstrAddr[9])
         );
  LHQD1BWP \nextInstrAddr_reg[10]  ( .E(N4162), .D(N4164), .Q(
        nextInstrAddr[10]) );
  LHQD1BWP \nextInstrAddr_reg[11]  ( .E(N4162), .D(N4165), .Q(
        nextInstrAddr[11]) );
  LHQD1BWP \nextInstrAddr_reg[12]  ( .E(N4162), .D(N4166), .Q(
        nextInstrAddr[12]) );
  LHQD1BWP \nextInstrAddr_reg[13]  ( .E(N4162), .D(N4167), .Q(
        nextInstrAddr[13]) );
  LHQD1BWP \nextInstrAddr_reg[14]  ( .E(N4162), .D(N4168), .Q(
        nextInstrAddr[14]) );
  LHQD1BWP \nextInstrAddr_reg[15]  ( .E(N4162), .D(N4169), .Q(
        nextInstrAddr[15]) );
  LHQD1BWP \nextInstrAddr_reg[8]  ( .E(N4162), .D(N4161), .Q(nextInstrAddr[8])
         );
  LHQD1BWP \nextInstrAddr_reg[7]  ( .E(N4162), .D(N4160), .Q(nextInstrAddr[7])
         );
  LHQD1BWP \nextInstrAddr_reg[6]  ( .E(N4162), .D(N4159), .Q(nextInstrAddr[6])
         );
  LHQD1BWP \nextInstrAddr_reg[5]  ( .E(N4162), .D(N4158), .Q(nextInstrAddr[5])
         );
  LHQD1BWP \nextInstrAddr_reg[4]  ( .E(N4162), .D(N4157), .Q(nextInstrAddr[4])
         );
  LHQD1BWP \nextInstrAddr_reg[3]  ( .E(N4162), .D(N4156), .Q(nextInstrAddr[3])
         );
  LHQD1BWP \nextInstrAddr_reg[2]  ( .E(N4162), .D(N4155), .Q(nextInstrAddr[2])
         );
  LHQD1BWP \nextInstrAddr_reg[1]  ( .E(N4162), .D(N4154), .Q(nextInstrAddr[1])
         );
  LHQD1BWP \nextInstrAddr_reg[0]  ( .E(N4162), .D(N4153), .Q(nextInstrAddr[0])
         );
  LHD4BWP \cycles_reg[0]  ( .E(N4170), .D(N4171), .Q(cycles[0]), .QN(n137) );
  LHD4BWP \cycles_reg[1]  ( .E(N4170), .D(N4172), .Q(cycles[1]), .QN(n136) );
  LHD4BWP \cycles_reg[2]  ( .E(N4170), .D(N4173), .Q(cycles[2]), .QN(n134) );
  LHD4BWP \cycles_reg[3]  ( .E(N4170), .D(N4174), .Q(cycles[3]), .QN(n132) );
  LHQD1BWP \cycles_reg[4]  ( .E(N4170), .D(N4175), .Q(cycles[4]) );
  LHQD1BWP \vectorToLoad_reg[255]  ( .E(n3582), .D(N4474), .Q(
        vectorToLoad[255]) );
  LHQD1BWP \vectorToLoad_reg[254]  ( .E(n3582), .D(N4473), .Q(
        vectorToLoad[254]) );
  LHQD1BWP \vectorToLoad_reg[253]  ( .E(n3582), .D(N4472), .Q(
        vectorToLoad[253]) );
  LHQD1BWP \vectorToLoad_reg[252]  ( .E(n3582), .D(N4471), .Q(
        vectorToLoad[252]) );
  LHQD1BWP \vectorToLoad_reg[251]  ( .E(n3582), .D(N4470), .Q(
        vectorToLoad[251]) );
  LHQD1BWP \vectorToLoad_reg[250]  ( .E(n3582), .D(N4469), .Q(
        vectorToLoad[250]) );
  LHQD1BWP \vectorToLoad_reg[249]  ( .E(n3582), .D(N4468), .Q(
        vectorToLoad[249]) );
  LHQD1BWP \vectorToLoad_reg[248]  ( .E(n3582), .D(N4467), .Q(
        vectorToLoad[248]) );
  LHQD1BWP \vectorToLoad_reg[247]  ( .E(n3600), .D(N4466), .Q(
        vectorToLoad[247]) );
  LHQD1BWP \vectorToLoad_reg[246]  ( .E(n3582), .D(N4465), .Q(
        vectorToLoad[246]) );
  LHQD1BWP \vectorToLoad_reg[245]  ( .E(n3600), .D(N4464), .Q(
        vectorToLoad[245]) );
  LHQD1BWP \vectorToLoad_reg[244]  ( .E(n3600), .D(N4463), .Q(
        vectorToLoad[244]) );
  LHQD1BWP \vectorToLoad_reg[243]  ( .E(n3582), .D(N4462), .Q(
        vectorToLoad[243]) );
  LHQD1BWP \vectorToLoad_reg[242]  ( .E(n3600), .D(N4461), .Q(
        vectorToLoad[242]) );
  LHQD1BWP \vectorToLoad_reg[241]  ( .E(n3582), .D(N4460), .Q(
        vectorToLoad[241]) );
  LHQD1BWP \vectorToLoad_reg[240]  ( .E(n3600), .D(N4459), .Q(
        vectorToLoad[240]) );
  LHQD1BWP \vectorToLoad_reg[239]  ( .E(n3582), .D(N4458), .Q(
        vectorToLoad[239]) );
  LHQD1BWP \vectorToLoad_reg[238]  ( .E(n3582), .D(N4457), .Q(
        vectorToLoad[238]) );
  LHQD1BWP \vectorToLoad_reg[237]  ( .E(n3582), .D(N4456), .Q(
        vectorToLoad[237]) );
  LHQD1BWP \vectorToLoad_reg[236]  ( .E(n3600), .D(N4455), .Q(
        vectorToLoad[236]) );
  LHQD1BWP \vectorToLoad_reg[235]  ( .E(n3582), .D(N4454), .Q(
        vectorToLoad[235]) );
  LHQD1BWP \vectorToLoad_reg[234]  ( .E(n3600), .D(N4453), .Q(
        vectorToLoad[234]) );
  LHQD1BWP \vectorToLoad_reg[233]  ( .E(n3582), .D(N4452), .Q(
        vectorToLoad[233]) );
  LHQD1BWP \vectorToLoad_reg[232]  ( .E(n3582), .D(N4451), .Q(
        vectorToLoad[232]) );
  LHQD1BWP \vectorToLoad_reg[231]  ( .E(n3582), .D(N4450), .Q(
        vectorToLoad[231]) );
  LHQD1BWP \vectorToLoad_reg[230]  ( .E(n3600), .D(N4449), .Q(
        vectorToLoad[230]) );
  LHQD1BWP \vectorToLoad_reg[229]  ( .E(n3582), .D(N4448), .Q(
        vectorToLoad[229]) );
  LHQD1BWP \vectorToLoad_reg[228]  ( .E(n3600), .D(N4447), .Q(
        vectorToLoad[228]) );
  LHQD1BWP \vectorToLoad_reg[227]  ( .E(n3600), .D(N4446), .Q(
        vectorToLoad[227]) );
  LHQD1BWP \vectorToLoad_reg[226]  ( .E(n3582), .D(N4445), .Q(
        vectorToLoad[226]) );
  LHQD1BWP \vectorToLoad_reg[225]  ( .E(n4630), .D(N4444), .Q(
        vectorToLoad[225]) );
  LHQD1BWP \vectorToLoad_reg[224]  ( .E(n3600), .D(N4443), .Q(
        vectorToLoad[224]) );
  LHQD1BWP \vectorToLoad_reg[223]  ( .E(n3600), .D(N4442), .Q(
        vectorToLoad[223]) );
  LHQD1BWP \vectorToLoad_reg[222]  ( .E(n3582), .D(N4441), .Q(
        vectorToLoad[222]) );
  LHQD1BWP \vectorToLoad_reg[221]  ( .E(n3600), .D(N4440), .Q(
        vectorToLoad[221]) );
  LHQD1BWP \vectorToLoad_reg[220]  ( .E(n3600), .D(N4439), .Q(
        vectorToLoad[220]) );
  LHQD1BWP \vectorToLoad_reg[219]  ( .E(n3582), .D(N4438), .Q(
        vectorToLoad[219]) );
  LHQD1BWP \vectorToLoad_reg[218]  ( .E(n3600), .D(N4437), .Q(
        vectorToLoad[218]) );
  LHQD1BWP \vectorToLoad_reg[217]  ( .E(n3582), .D(N4436), .Q(
        vectorToLoad[217]) );
  LHQD1BWP \vectorToLoad_reg[216]  ( .E(n3582), .D(N4435), .Q(
        vectorToLoad[216]) );
  LHQD1BWP \vectorToLoad_reg[215]  ( .E(n3600), .D(N4434), .Q(
        vectorToLoad[215]) );
  LHQD1BWP \vectorToLoad_reg[214]  ( .E(n3582), .D(N4433), .Q(
        vectorToLoad[214]) );
  LHQD1BWP \vectorToLoad_reg[213]  ( .E(n3600), .D(N4431), .Q(
        vectorToLoad[213]) );
  LHQD1BWP \vectorToLoad_reg[212]  ( .E(n3600), .D(N4430), .Q(
        vectorToLoad[212]) );
  LHQD1BWP \vectorToLoad_reg[211]  ( .E(n3600), .D(N4429), .Q(
        vectorToLoad[211]) );
  LHQD1BWP \vectorToLoad_reg[210]  ( .E(n4630), .D(N4428), .Q(
        vectorToLoad[210]) );
  LHQD1BWP \vectorToLoad_reg[209]  ( .E(n3582), .D(N4427), .Q(
        vectorToLoad[209]) );
  LHQD1BWP \vectorToLoad_reg[208]  ( .E(n3582), .D(N4426), .Q(
        vectorToLoad[208]) );
  LHQD1BWP \vectorToLoad_reg[207]  ( .E(n3600), .D(N4425), .Q(
        vectorToLoad[207]) );
  LHQD1BWP \vectorToLoad_reg[206]  ( .E(n3582), .D(N4424), .Q(
        vectorToLoad[206]) );
  LHQD1BWP \vectorToLoad_reg[205]  ( .E(n3582), .D(N4423), .Q(
        vectorToLoad[205]) );
  LHQD1BWP \vectorToLoad_reg[204]  ( .E(n3582), .D(N4422), .Q(
        vectorToLoad[204]) );
  LHQD1BWP \vectorToLoad_reg[203]  ( .E(n3582), .D(N4421), .Q(
        vectorToLoad[203]) );
  LHQD1BWP \vectorToLoad_reg[202]  ( .E(n3582), .D(N4420), .Q(
        vectorToLoad[202]) );
  LHQD1BWP \vectorToLoad_reg[201]  ( .E(n4630), .D(N4419), .Q(
        vectorToLoad[201]) );
  LHQD1BWP \vectorToLoad_reg[200]  ( .E(n3600), .D(N4418), .Q(
        vectorToLoad[200]) );
  LHQD1BWP \vectorToLoad_reg[199]  ( .E(n3600), .D(N4417), .Q(
        vectorToLoad[199]) );
  LHQD1BWP \vectorToLoad_reg[198]  ( .E(n3582), .D(N4416), .Q(
        vectorToLoad[198]) );
  LHQD1BWP \vectorToLoad_reg[197]  ( .E(n3582), .D(N4415), .Q(
        vectorToLoad[197]) );
  LHQD1BWP \vectorToLoad_reg[196]  ( .E(n3600), .D(N4414), .Q(
        vectorToLoad[196]) );
  LHQD1BWP \vectorToLoad_reg[195]  ( .E(n3600), .D(N4413), .Q(
        vectorToLoad[195]) );
  LHQD1BWP \vectorToLoad_reg[194]  ( .E(n3582), .D(N4412), .Q(
        vectorToLoad[194]) );
  LHQD1BWP \vectorToLoad_reg[193]  ( .E(n3600), .D(N4411), .Q(
        vectorToLoad[193]) );
  LHQD1BWP \vectorToLoad_reg[192]  ( .E(n3600), .D(N4410), .Q(
        vectorToLoad[192]) );
  LHQD1BWP \vectorToLoad_reg[191]  ( .E(n3582), .D(N4409), .Q(
        vectorToLoad[191]) );
  LHQD1BWP \vectorToLoad_reg[190]  ( .E(n3600), .D(N4408), .Q(
        vectorToLoad[190]) );
  LHQD1BWP \vectorToLoad_reg[189]  ( .E(n3582), .D(N4407), .Q(
        vectorToLoad[189]) );
  LHQD1BWP \vectorToLoad_reg[188]  ( .E(n3600), .D(N4406), .Q(
        vectorToLoad[188]) );
  LHQD1BWP \vectorToLoad_reg[187]  ( .E(n3582), .D(N4405), .Q(
        vectorToLoad[187]) );
  LHQD1BWP \vectorToLoad_reg[186]  ( .E(n3600), .D(N4404), .Q(
        vectorToLoad[186]) );
  LHQD1BWP \vectorToLoad_reg[185]  ( .E(n3582), .D(N4403), .Q(
        vectorToLoad[185]) );
  LHQD1BWP \vectorToLoad_reg[184]  ( .E(n4630), .D(N4402), .Q(
        vectorToLoad[184]) );
  LHQD1BWP \vectorToLoad_reg[183]  ( .E(n4630), .D(N4401), .Q(
        vectorToLoad[183]) );
  LHQD1BWP \vectorToLoad_reg[182]  ( .E(n3600), .D(N4400), .Q(
        vectorToLoad[182]) );
  LHQD1BWP \vectorToLoad_reg[181]  ( .E(n3600), .D(N4399), .Q(
        vectorToLoad[181]) );
  LHQD1BWP \vectorToLoad_reg[180]  ( .E(n3582), .D(N4398), .Q(
        vectorToLoad[180]) );
  LHQD1BWP \vectorToLoad_reg[179]  ( .E(n3600), .D(N4397), .Q(
        vectorToLoad[179]) );
  LHQD1BWP \vectorToLoad_reg[178]  ( .E(n3600), .D(N4396), .Q(
        vectorToLoad[178]) );
  LHQD1BWP \vectorToLoad_reg[177]  ( .E(n3582), .D(N4395), .Q(
        vectorToLoad[177]) );
  LHQD1BWP \vectorToLoad_reg[176]  ( .E(n3600), .D(N4394), .Q(
        vectorToLoad[176]) );
  LHQD1BWP \vectorToLoad_reg[175]  ( .E(n3600), .D(N4393), .Q(
        vectorToLoad[175]) );
  LHQD1BWP \vectorToLoad_reg[174]  ( .E(n3582), .D(N4392), .Q(
        vectorToLoad[174]) );
  LHQD1BWP \vectorToLoad_reg[173]  ( .E(n3582), .D(N4391), .Q(
        vectorToLoad[173]) );
  LHQD1BWP \vectorToLoad_reg[172]  ( .E(n4630), .D(N4390), .Q(
        vectorToLoad[172]) );
  LHQD1BWP \vectorToLoad_reg[171]  ( .E(n4630), .D(N4389), .Q(
        vectorToLoad[171]) );
  LHQD1BWP \vectorToLoad_reg[170]  ( .E(n4630), .D(N4388), .Q(
        vectorToLoad[170]) );
  LHQD1BWP \vectorToLoad_reg[169]  ( .E(n3600), .D(N4387), .Q(
        vectorToLoad[169]) );
  LHQD1BWP \vectorToLoad_reg[168]  ( .E(n3582), .D(N4386), .Q(
        vectorToLoad[168]) );
  LHQD1BWP \vectorToLoad_reg[167]  ( .E(n3600), .D(N4385), .Q(
        vectorToLoad[167]) );
  LHQD1BWP \vectorToLoad_reg[166]  ( .E(n4630), .D(N4384), .Q(
        vectorToLoad[166]) );
  LHQD1BWP \vectorToLoad_reg[165]  ( .E(n4630), .D(N4383), .Q(
        vectorToLoad[165]) );
  LHQD1BWP \vectorToLoad_reg[164]  ( .E(n3600), .D(N4382), .Q(
        vectorToLoad[164]) );
  LHQD1BWP \vectorToLoad_reg[163]  ( .E(n3600), .D(N4381), .Q(
        vectorToLoad[163]) );
  LHQD1BWP \vectorToLoad_reg[162]  ( .E(n3582), .D(N4380), .Q(
        vectorToLoad[162]) );
  LHQD1BWP \vectorToLoad_reg[161]  ( .E(n4630), .D(N4379), .Q(
        vectorToLoad[161]) );
  LHQD1BWP \vectorToLoad_reg[160]  ( .E(n4630), .D(N4378), .Q(
        vectorToLoad[160]) );
  LHQD1BWP \vectorToLoad_reg[159]  ( .E(n4630), .D(N4377), .Q(
        vectorToLoad[159]) );
  LHQD1BWP \vectorToLoad_reg[158]  ( .E(n3600), .D(N4376), .Q(
        vectorToLoad[158]) );
  LHQD1BWP \vectorToLoad_reg[157]  ( .E(n3600), .D(N4375), .Q(
        vectorToLoad[157]) );
  LHQD1BWP \vectorToLoad_reg[156]  ( .E(n3582), .D(N4374), .Q(
        vectorToLoad[156]) );
  LHQD1BWP \vectorToLoad_reg[155]  ( .E(n4630), .D(N4373), .Q(
        vectorToLoad[155]) );
  LHQD1BWP \vectorToLoad_reg[154]  ( .E(n3600), .D(N4372), .Q(
        vectorToLoad[154]) );
  LHQD1BWP \vectorToLoad_reg[153]  ( .E(n3582), .D(N4371), .Q(
        vectorToLoad[153]) );
  LHQD1BWP \vectorToLoad_reg[152]  ( .E(n3582), .D(N4370), .Q(
        vectorToLoad[152]) );
  LHQD1BWP \vectorToLoad_reg[151]  ( .E(n4630), .D(N4369), .Q(
        vectorToLoad[151]) );
  LHQD1BWP \vectorToLoad_reg[150]  ( .E(n4630), .D(N4368), .Q(
        vectorToLoad[150]) );
  LHQD1BWP \vectorToLoad_reg[149]  ( .E(n3582), .D(N4367), .Q(
        vectorToLoad[149]) );
  LHQD1BWP \vectorToLoad_reg[148]  ( .E(n3582), .D(N4366), .Q(
        vectorToLoad[148]) );
  LHQD1BWP \vectorToLoad_reg[147]  ( .E(n3600), .D(N4365), .Q(
        vectorToLoad[147]) );
  LHQD1BWP \vectorToLoad_reg[146]  ( .E(n4630), .D(N4364), .Q(
        vectorToLoad[146]) );
  LHQD1BWP \vectorToLoad_reg[145]  ( .E(n3600), .D(N4363), .Q(
        vectorToLoad[145]) );
  LHQD1BWP \vectorToLoad_reg[144]  ( .E(n3600), .D(N4362), .Q(
        vectorToLoad[144]) );
  LHQD1BWP \vectorToLoad_reg[143]  ( .E(n3600), .D(N4361), .Q(
        vectorToLoad[143]) );
  LHQD1BWP \vectorToLoad_reg[142]  ( .E(n3600), .D(N4360), .Q(
        vectorToLoad[142]) );
  LHQD1BWP \vectorToLoad_reg[141]  ( .E(n3582), .D(N4359), .Q(
        vectorToLoad[141]) );
  LHQD1BWP \vectorToLoad_reg[140]  ( .E(n3600), .D(N4358), .Q(
        vectorToLoad[140]) );
  LHQD1BWP \vectorToLoad_reg[139]  ( .E(n4630), .D(N4357), .Q(
        vectorToLoad[139]) );
  LHQD1BWP \vectorToLoad_reg[138]  ( .E(n3582), .D(N4356), .Q(
        vectorToLoad[138]) );
  LHQD1BWP \vectorToLoad_reg[137]  ( .E(n3582), .D(N4355), .Q(
        vectorToLoad[137]) );
  LHQD1BWP \vectorToLoad_reg[136]  ( .E(n3582), .D(N4354), .Q(
        vectorToLoad[136]) );
  LHQD1BWP \vectorToLoad_reg[135]  ( .E(n3582), .D(N4353), .Q(
        vectorToLoad[135]) );
  LHQD1BWP \vectorToLoad_reg[134]  ( .E(n3582), .D(N4352), .Q(
        vectorToLoad[134]) );
  LHQD1BWP \vectorToLoad_reg[133]  ( .E(n3582), .D(N4351), .Q(
        vectorToLoad[133]) );
  LHQD1BWP \vectorToLoad_reg[132]  ( .E(n3600), .D(N4350), .Q(
        vectorToLoad[132]) );
  LHQD1BWP \vectorToLoad_reg[131]  ( .E(n3582), .D(N4349), .Q(
        vectorToLoad[131]) );
  LHQD1BWP \vectorToLoad_reg[130]  ( .E(n3600), .D(N4348), .Q(
        vectorToLoad[130]) );
  LHQD1BWP \vectorToLoad_reg[129]  ( .E(n3600), .D(N4347), .Q(
        vectorToLoad[129]) );
  LHQD1BWP \vectorToLoad_reg[128]  ( .E(n4630), .D(N4346), .Q(
        vectorToLoad[128]) );
  LHQD1BWP \vectorToLoad_reg[99]  ( .E(n3582), .D(N4316), .Q(vectorToLoad[99])
         );
  LHQD1BWP \vectorToLoad_reg[98]  ( .E(n3600), .D(N4315), .Q(vectorToLoad[98])
         );
  LHQD1BWP \vectorToLoad_reg[97]  ( .E(n3582), .D(N4314), .Q(vectorToLoad[97])
         );
  LHQD1BWP \vectorToLoad_reg[96]  ( .E(n3600), .D(N4313), .Q(vectorToLoad[96])
         );
  LHQD1BWP \vectorToLoad_reg[95]  ( .E(n3582), .D(N4312), .Q(vectorToLoad[95])
         );
  LHQD1BWP \vectorToLoad_reg[94]  ( .E(n3600), .D(N4311), .Q(vectorToLoad[94])
         );
  LHQD1BWP \vectorToLoad_reg[93]  ( .E(n3582), .D(N4310), .Q(vectorToLoad[93])
         );
  LHQD1BWP \vectorToLoad_reg[92]  ( .E(n3600), .D(N4309), .Q(vectorToLoad[92])
         );
  LHQD1BWP \vectorToLoad_reg[91]  ( .E(n3600), .D(N4308), .Q(vectorToLoad[91])
         );
  LHQD1BWP \vectorToLoad_reg[90]  ( .E(n3582), .D(N4307), .Q(vectorToLoad[90])
         );
  LHQD1BWP \vectorToLoad_reg[89]  ( .E(n3600), .D(N4306), .Q(vectorToLoad[89])
         );
  LHQD1BWP \vectorToLoad_reg[88]  ( .E(n3582), .D(N4305), .Q(vectorToLoad[88])
         );
  LHQD1BWP \vectorToLoad_reg[87]  ( .E(n3600), .D(N4304), .Q(vectorToLoad[87])
         );
  LHQD1BWP \vectorToLoad_reg[86]  ( .E(n3582), .D(N4303), .Q(vectorToLoad[86])
         );
  LHQD1BWP \vectorToLoad_reg[85]  ( .E(n3600), .D(N4302), .Q(vectorToLoad[85])
         );
  LHQD1BWP \vectorToLoad_reg[84]  ( .E(n3582), .D(N4301), .Q(vectorToLoad[84])
         );
  LHQD1BWP \vectorToLoad_reg[83]  ( .E(n3582), .D(N4300), .Q(vectorToLoad[83])
         );
  LHQD1BWP \vectorToLoad_reg[82]  ( .E(n3582), .D(N4299), .Q(vectorToLoad[82])
         );
  LHQD1BWP \vectorToLoad_reg[81]  ( .E(n3600), .D(N4298), .Q(vectorToLoad[81])
         );
  LHQD1BWP \vectorToLoad_reg[80]  ( .E(n3600), .D(N4297), .Q(vectorToLoad[80])
         );
  LHQD1BWP \vectorToLoad_reg[79]  ( .E(n3600), .D(N4296), .Q(vectorToLoad[79])
         );
  LHQD1BWP \vectorToLoad_reg[78]  ( .E(n3600), .D(N4295), .Q(vectorToLoad[78])
         );
  LHQD1BWP \vectorToLoad_reg[77]  ( .E(n3600), .D(N4294), .Q(vectorToLoad[77])
         );
  LHQD1BWP \vectorToLoad_reg[76]  ( .E(n3600), .D(N4293), .Q(vectorToLoad[76])
         );
  LHQD1BWP \vectorToLoad_reg[75]  ( .E(n3600), .D(N4292), .Q(vectorToLoad[75])
         );
  LHQD1BWP \vectorToLoad_reg[74]  ( .E(n3600), .D(N4291), .Q(vectorToLoad[74])
         );
  LHQD1BWP \vectorToLoad_reg[73]  ( .E(n3600), .D(N4290), .Q(vectorToLoad[73])
         );
  LHQD1BWP \vectorToLoad_reg[72]  ( .E(n3600), .D(N4289), .Q(vectorToLoad[72])
         );
  LHQD1BWP \vectorToLoad_reg[71]  ( .E(n3600), .D(N4288), .Q(vectorToLoad[71])
         );
  LHQD1BWP \vectorToLoad_reg[70]  ( .E(n3600), .D(N4287), .Q(vectorToLoad[70])
         );
  LHQD1BWP \vectorToLoad_reg[69]  ( .E(n3582), .D(N4286), .Q(vectorToLoad[69])
         );
  LHQD1BWP \vectorToLoad_reg[68]  ( .E(n3582), .D(N4285), .Q(vectorToLoad[68])
         );
  LHQD1BWP \vectorToLoad_reg[67]  ( .E(n3582), .D(N4284), .Q(vectorToLoad[67])
         );
  LHQD1BWP \vectorToLoad_reg[66]  ( .E(n3582), .D(N4283), .Q(vectorToLoad[66])
         );
  LHQD1BWP \vectorToLoad_reg[65]  ( .E(n3582), .D(N4282), .Q(vectorToLoad[65])
         );
  LHQD1BWP \vectorToLoad_reg[64]  ( .E(n3582), .D(N4281), .Q(vectorToLoad[64])
         );
  LHQD1BWP \vectorToLoad_reg[63]  ( .E(n3582), .D(N4280), .Q(vectorToLoad[63])
         );
  LHQD1BWP \vectorToLoad_reg[62]  ( .E(n3582), .D(N4279), .Q(vectorToLoad[62])
         );
  LHQD1BWP \vectorToLoad_reg[61]  ( .E(n3582), .D(N4278), .Q(vectorToLoad[61])
         );
  LHQD1BWP \vectorToLoad_reg[60]  ( .E(n3582), .D(N4277), .Q(vectorToLoad[60])
         );
  LHQD1BWP \vectorToLoad_reg[59]  ( .E(n3582), .D(N4276), .Q(vectorToLoad[59])
         );
  LHQD1BWP \vectorToLoad_reg[58]  ( .E(n3582), .D(N4275), .Q(vectorToLoad[58])
         );
  LHQD1BWP \vectorToLoad_reg[57]  ( .E(n3600), .D(N4274), .Q(vectorToLoad[57])
         );
  LHQD1BWP \vectorToLoad_reg[56]  ( .E(n3600), .D(N4273), .Q(vectorToLoad[56])
         );
  LHQD1BWP \vectorToLoad_reg[55]  ( .E(n3600), .D(N4272), .Q(vectorToLoad[55])
         );
  LHQD1BWP \vectorToLoad_reg[54]  ( .E(n3600), .D(N4271), .Q(vectorToLoad[54])
         );
  LHQD1BWP \vectorToLoad_reg[53]  ( .E(n3600), .D(N4270), .Q(vectorToLoad[53])
         );
  LHQD1BWP \vectorToLoad_reg[52]  ( .E(n3600), .D(N4269), .Q(vectorToLoad[52])
         );
  LHQD1BWP \vectorToLoad_reg[51]  ( .E(n3600), .D(N4268), .Q(vectorToLoad[51])
         );
  LHQD1BWP \vectorToLoad_reg[50]  ( .E(n3600), .D(N4267), .Q(vectorToLoad[50])
         );
  LHQD1BWP \vectorToLoad_reg[49]  ( .E(n3600), .D(N4266), .Q(vectorToLoad[49])
         );
  LHQD1BWP \vectorToLoad_reg[48]  ( .E(n3600), .D(N4265), .Q(vectorToLoad[48])
         );
  LHQD1BWP \vectorToLoad_reg[47]  ( .E(n3600), .D(N4264), .Q(vectorToLoad[47])
         );
  LHQD1BWP \vectorToLoad_reg[46]  ( .E(n3600), .D(N4263), .Q(vectorToLoad[46])
         );
  LHQD1BWP \vectorToLoad_reg[45]  ( .E(n3600), .D(N4262), .Q(vectorToLoad[45])
         );
  LHQD1BWP \vectorToLoad_reg[44]  ( .E(n3582), .D(N4261), .Q(vectorToLoad[44])
         );
  LHQD1BWP \vectorToLoad_reg[43]  ( .E(n3600), .D(N4260), .Q(vectorToLoad[43])
         );
  LHQD1BWP \vectorToLoad_reg[42]  ( .E(n3582), .D(N4259), .Q(vectorToLoad[42])
         );
  LHQD1BWP \vectorToLoad_reg[41]  ( .E(n3600), .D(N4258), .Q(vectorToLoad[41])
         );
  LHQD1BWP \vectorToLoad_reg[40]  ( .E(n3582), .D(N4257), .Q(vectorToLoad[40])
         );
  LHQD1BWP \vectorToLoad_reg[39]  ( .E(n3600), .D(N4256), .Q(vectorToLoad[39])
         );
  LHQD1BWP \vectorToLoad_reg[38]  ( .E(n3582), .D(N4255), .Q(vectorToLoad[38])
         );
  LHQD1BWP \vectorToLoad_reg[37]  ( .E(n3600), .D(N4254), .Q(vectorToLoad[37])
         );
  LHQD1BWP \vectorToLoad_reg[36]  ( .E(n3582), .D(N4253), .Q(vectorToLoad[36])
         );
  LHQD1BWP \vectorToLoad_reg[35]  ( .E(n3600), .D(N4252), .Q(vectorToLoad[35])
         );
  LHQD1BWP \vectorToLoad_reg[34]  ( .E(n3582), .D(N4251), .Q(vectorToLoad[34])
         );
  LHQD1BWP \vectorToLoad_reg[33]  ( .E(n3582), .D(N4250), .Q(vectorToLoad[33])
         );
  LHQD1BWP \vectorToLoad_reg[32]  ( .E(n3582), .D(N4249), .Q(vectorToLoad[32])
         );
  LHQD1BWP \vectorToLoad_reg[31]  ( .E(n3582), .D(N4248), .Q(vectorToLoad[31])
         );
  LHQD1BWP \vectorToLoad_reg[30]  ( .E(n3600), .D(N4247), .Q(vectorToLoad[30])
         );
  LHQD1BWP \vectorToLoad_reg[29]  ( .E(n3582), .D(N4246), .Q(vectorToLoad[29])
         );
  LHQD1BWP \vectorToLoad_reg[28]  ( .E(n3600), .D(N4245), .Q(vectorToLoad[28])
         );
  LHQD1BWP \vectorToLoad_reg[27]  ( .E(n3582), .D(N4244), .Q(vectorToLoad[27])
         );
  LHQD1BWP \vectorToLoad_reg[26]  ( .E(n4630), .D(N4243), .Q(vectorToLoad[26])
         );
  LHQD1BWP \vectorToLoad_reg[25]  ( .E(n3582), .D(N4242), .Q(vectorToLoad[25])
         );
  LHQD1BWP \vectorToLoad_reg[24]  ( .E(n4630), .D(N4241), .Q(vectorToLoad[24])
         );
  LHQD1BWP \vectorToLoad_reg[23]  ( .E(n4630), .D(N4240), .Q(vectorToLoad[23])
         );
  LHQD1BWP \vectorToLoad_reg[22]  ( .E(n4630), .D(N4239), .Q(vectorToLoad[22])
         );
  LHQD1BWP \vectorToLoad_reg[21]  ( .E(n4630), .D(N4238), .Q(vectorToLoad[21])
         );
  LHQD1BWP \vectorToLoad_reg[20]  ( .E(n3582), .D(N4237), .Q(vectorToLoad[20])
         );
  LHQD1BWP \vectorToLoad_reg[19]  ( .E(n3582), .D(N4236), .Q(vectorToLoad[19])
         );
  LHQD1BWP \vectorToLoad_reg[18]  ( .E(n3600), .D(N4235), .Q(vectorToLoad[18])
         );
  LHQD1BWP \vectorToLoad_reg[17]  ( .E(n3582), .D(N4234), .Q(vectorToLoad[17])
         );
  LHQD1BWP \vectorToLoad_reg[16]  ( .E(n3582), .D(N4233), .Q(vectorToLoad[16])
         );
  LHQD1BWP \vectorToLoad_reg[127]  ( .E(n3600), .D(N4345), .Q(
        vectorToLoad[127]) );
  LHQD1BWP \vectorToLoad_reg[126]  ( .E(n3600), .D(N4344), .Q(
        vectorToLoad[126]) );
  LHQD1BWP \vectorToLoad_reg[125]  ( .E(n3600), .D(N4343), .Q(
        vectorToLoad[125]) );
  LHQD1BWP \vectorToLoad_reg[124]  ( .E(n3600), .D(N4342), .Q(
        vectorToLoad[124]) );
  LHQD1BWP \vectorToLoad_reg[123]  ( .E(n3582), .D(N4341), .Q(
        vectorToLoad[123]) );
  LHQD1BWP \vectorToLoad_reg[122]  ( .E(n3582), .D(N4340), .Q(
        vectorToLoad[122]) );
  LHQD1BWP \vectorToLoad_reg[121]  ( .E(n3600), .D(N4339), .Q(
        vectorToLoad[121]) );
  LHQD1BWP \vectorToLoad_reg[120]  ( .E(n4630), .D(N4338), .Q(
        vectorToLoad[120]) );
  LHQD1BWP \vectorToLoad_reg[119]  ( .E(n3600), .D(N4337), .Q(
        vectorToLoad[119]) );
  LHQD1BWP \vectorToLoad_reg[118]  ( .E(n3582), .D(N4336), .Q(
        vectorToLoad[118]) );
  LHQD1BWP \vectorToLoad_reg[117]  ( .E(n3600), .D(N4335), .Q(
        vectorToLoad[117]) );
  LHQD1BWP \vectorToLoad_reg[116]  ( .E(n3582), .D(N4334), .Q(
        vectorToLoad[116]) );
  LHQD1BWP \vectorToLoad_reg[115]  ( .E(n3600), .D(N4333), .Q(
        vectorToLoad[115]) );
  LHQD1BWP \vectorToLoad_reg[114]  ( .E(n3582), .D(N4331), .Q(
        vectorToLoad[114]) );
  LHQD1BWP \vectorToLoad_reg[113]  ( .E(n3600), .D(N4330), .Q(
        vectorToLoad[113]) );
  LHQD1BWP \vectorToLoad_reg[112]  ( .E(n3582), .D(N4329), .Q(
        vectorToLoad[112]) );
  LHQD1BWP \vectorToLoad_reg[111]  ( .E(n3600), .D(N4328), .Q(
        vectorToLoad[111]) );
  LHQD1BWP \vectorToLoad_reg[110]  ( .E(n3582), .D(N4327), .Q(
        vectorToLoad[110]) );
  LHQD1BWP \vectorToLoad_reg[109]  ( .E(n3600), .D(N4326), .Q(
        vectorToLoad[109]) );
  LHQD1BWP \vectorToLoad_reg[108]  ( .E(n3582), .D(N4325), .Q(
        vectorToLoad[108]) );
  LHQD1BWP \vectorToLoad_reg[107]  ( .E(n3600), .D(N4324), .Q(
        vectorToLoad[107]) );
  LHQD1BWP \vectorToLoad_reg[106]  ( .E(n3582), .D(N4323), .Q(
        vectorToLoad[106]) );
  LHQD1BWP \vectorToLoad_reg[105]  ( .E(n3600), .D(N4322), .Q(
        vectorToLoad[105]) );
  LHQD1BWP \vectorToLoad_reg[104]  ( .E(n3600), .D(N4321), .Q(
        vectorToLoad[104]) );
  LHQD1BWP \vectorToLoad_reg[103]  ( .E(n3582), .D(N4320), .Q(
        vectorToLoad[103]) );
  LHQD1BWP \vectorToLoad_reg[102]  ( .E(n3600), .D(N4319), .Q(
        vectorToLoad[102]) );
  LHQD1BWP \vectorToLoad_reg[101]  ( .E(n3582), .D(N4318), .Q(
        vectorToLoad[101]) );
  LHQD1BWP \vectorToLoad_reg[100]  ( .E(n3582), .D(N4317), .Q(
        vectorToLoad[100]) );
  LHQD1BWP \memAddr_reg[0]  ( .E(N4133), .D(N4134), .Q(Addr[0]) );
  LHQD1BWP \memAddr_reg[1]  ( .E(N4133), .D(N4135), .Q(Addr[1]) );
  LHQD1BWP \memAddr_reg[2]  ( .E(N4133), .D(N4136), .Q(Addr[2]) );
  LHQD1BWP \memAddr_reg[3]  ( .E(N4133), .D(N4137), .Q(Addr[3]) );
  LHQD1BWP \memAddr_reg[4]  ( .E(N4133), .D(N4138), .Q(Addr[4]) );
  LHQD1BWP \memAddr_reg[5]  ( .E(N4133), .D(N4139), .Q(Addr[5]) );
  LHQD1BWP \memAddr_reg[6]  ( .E(N4133), .D(N4140), .Q(Addr[6]) );
  LHQD1BWP \memAddr_reg[7]  ( .E(N4133), .D(N4141), .Q(Addr[7]) );
  LHQD1BWP \memAddr_reg[8]  ( .E(N4133), .D(N4142), .Q(Addr[8]) );
  LHQD1BWP \memAddr_reg[9]  ( .E(N4133), .D(N4143), .Q(Addr[9]) );
  LHQD1BWP \memAddr_reg[10]  ( .E(N4133), .D(N4144), .Q(Addr[10]) );
  LHQD1BWP \memAddr_reg[11]  ( .E(N4133), .D(N4145), .Q(Addr[11]) );
  LHQD1BWP \memAddr_reg[12]  ( .E(N4133), .D(N4146), .Q(Addr[12]) );
  LHQD1BWP \memAddr_reg[13]  ( .E(N4133), .D(N4147), .Q(Addr[13]) );
  LHQD1BWP \memAddr_reg[14]  ( .E(N4133), .D(N4148), .Q(Addr[14]) );
  LHQD1BWP \memAddr_reg[15]  ( .E(N4133), .D(N4149), .Q(Addr[15]) );
  LNQD1BWP \instrIn_reg[11]  ( .D(DataIn[11]), .EN(n3020), .Q(instrIn[11]) );
  LNQD1BWP \instrIn_reg[10]  ( .D(DataIn[10]), .EN(n3020), .Q(instrIn[10]) );
  LNQD1BWP \instrIn_reg[9]  ( .D(DataIn[9]), .EN(n3020), .Q(instrIn[9]) );
  LNQD1BWP \instrIn_reg[8]  ( .D(DataIn[8]), .EN(n3020), .Q(instrIn[8]) );
  LNQD1BWP \instrIn_reg[7]  ( .D(DataIn[7]), .EN(n3020), .Q(instrIn[7]) );
  LNQD1BWP \instrIn_reg[6]  ( .D(DataIn[6]), .EN(n3020), .Q(instrIn[6]) );
  LHQD1BWP \op2_reg[14]  ( .E(N4208), .D(N4206), .Q(\alu/N684 ) );
  LHQD1BWP \op2_reg[12]  ( .E(N4208), .D(N4204), .Q(op2[12]) );
  LHQD1BWP \op2_reg[11]  ( .E(N4208), .D(N4203), .Q(op2[11]) );
  LHQD1BWP \op2_reg[10]  ( .E(N4208), .D(N4202), .Q(op2[10]) );
  LNQD1BWP \instrIn_reg[4]  ( .D(DataIn[4]), .EN(n3020), .Q(instrIn[4]) );
  LHQD1BWP \op2_reg[4]  ( .E(N4208), .D(N4196), .Q(op2[4]) );
  LNQD1BWP \instrIn_reg[3]  ( .D(DataIn[3]), .EN(n3020), .Q(instrIn[3]) );
  LHQD1BWP \op2_reg[3]  ( .E(N4208), .D(N4195), .Q(op2[3]) );
  LNQD1BWP \instrIn_reg[2]  ( .D(DataIn[2]), .EN(n3020), .Q(instrIn[2]) );
  LHQD1BWP \op2_reg[2]  ( .E(N4208), .D(N4194), .Q(op2[2]) );
  LNQD1BWP \instrIn_reg[1]  ( .D(DataIn[1]), .EN(n3020), .Q(instrIn[1]) );
  LHQD1BWP \op2_reg[1]  ( .E(N4208), .D(N4193), .Q(op2[1]) );
  LNQD1BWP \instrIn_reg[0]  ( .D(DataIn[0]), .EN(n3020), .Q(instrIn[0]) );
  LHQD1BWP \op2_reg[0]  ( .E(N4208), .D(N4192), .Q(op2[0]) );
  LHQD1BWP \op1_reg[15]  ( .E(N4208), .D(N4191), .Q(op1[15]) );
  LHQD1BWP \op1_reg[14]  ( .E(N4208), .D(N4190), .Q(\alu/N683 ) );
  LHQD1BWP \op1_reg[12]  ( .E(N4208), .D(N4188), .Q(op1[12]) );
  LHQD1BWP \op1_reg[11]  ( .E(N4208), .D(N4187), .Q(op1[11]) );
  LHQD1BWP \op1_reg[10]  ( .E(N4208), .D(N4186), .Q(op1[10]) );
  LHQD1BWP \op1_reg[9]  ( .E(N4208), .D(N4185), .Q(op1[9]) );
  LHQD1BWP \op1_reg[8]  ( .E(N4208), .D(N4184), .Q(op1[8]) );
  LHQD1BWP \op1_reg[7]  ( .E(N4208), .D(N4183), .Q(op1[7]) );
  LHQD1BWP \op1_reg[6]  ( .E(N4208), .D(N4182), .Q(op1[6]) );
  LHQD1BWP \op1_reg[5]  ( .E(N4208), .D(N4181), .Q(op1[5]) );
  LHQD1BWP \op1_reg[4]  ( .E(N4208), .D(N4180), .Q(op1[4]) );
  LHQD1BWP \op1_reg[3]  ( .E(N4208), .D(N4179), .Q(op1[3]) );
  LHQD1BWP \op1_reg[2]  ( .E(N4208), .D(N4178), .Q(op1[2]) );
  LHQD1BWP \op1_reg[1]  ( .E(N4208), .D(N4177), .Q(op1[1]) );
  LHQD1BWP \op1_reg[0]  ( .E(N4208), .D(N4176), .Q(op1[0]) );
  LHQD1BWP overflow_reg ( .E(N4209), .D(N4210), .Q(overflow) );
  LHQD1BWP \vrf/regTable_reg[7][0]  ( .E(n3583), .D(\vrf/N18 ), .Q(
        \vrf/regTable[7][0] ) );
  LHQD1BWP \vrf/regTable_reg[7][1]  ( .E(n3583), .D(\vrf/N19 ), .Q(
        \vrf/regTable[7][1] ) );
  LHQD1BWP \vrf/regTable_reg[7][2]  ( .E(n3583), .D(\vrf/N20 ), .Q(
        \vrf/regTable[7][2] ) );
  LHQD1BWP \vrf/regTable_reg[7][3]  ( .E(n3583), .D(\vrf/N21 ), .Q(
        \vrf/regTable[7][3] ) );
  LHQD1BWP \vrf/regTable_reg[7][4]  ( .E(n3583), .D(\vrf/N22 ), .Q(
        \vrf/regTable[7][4] ) );
  LHQD1BWP \vrf/regTable_reg[7][5]  ( .E(n3583), .D(\vrf/N23 ), .Q(
        \vrf/regTable[7][5] ) );
  LHQD1BWP \vrf/regTable_reg[7][6]  ( .E(n3583), .D(\vrf/N24 ), .Q(
        \vrf/regTable[7][6] ) );
  LHQD1BWP \vrf/regTable_reg[7][7]  ( .E(n3583), .D(\vrf/N25 ), .Q(
        \vrf/regTable[7][7] ) );
  LHQD1BWP \vrf/regTable_reg[7][8]  ( .E(n3583), .D(\vrf/N26 ), .Q(
        \vrf/regTable[7][8] ) );
  LHQD1BWP \vrf/regTable_reg[7][9]  ( .E(n3583), .D(\vrf/N27 ), .Q(
        \vrf/regTable[7][9] ) );
  LHQD1BWP \vrf/regTable_reg[7][10]  ( .E(n3583), .D(\vrf/N28 ), .Q(
        \vrf/regTable[7][10] ) );
  LHQD1BWP \vrf/regTable_reg[7][11]  ( .E(n3583), .D(\vrf/N29 ), .Q(
        \vrf/regTable[7][11] ) );
  LHQD1BWP \vrf/regTable_reg[7][12]  ( .E(n3583), .D(\vrf/N30 ), .Q(
        \vrf/regTable[7][12] ) );
  LHQD1BWP \vrf/regTable_reg[7][13]  ( .E(n3583), .D(\vrf/N31 ), .Q(
        \vrf/regTable[7][13] ) );
  LHQD1BWP \vrf/regTable_reg[7][14]  ( .E(n3583), .D(\vrf/N32 ), .Q(
        \vrf/regTable[7][14] ) );
  LHQD1BWP \vrf/regTable_reg[7][15]  ( .E(n3583), .D(\vrf/N33 ), .Q(
        \vrf/regTable[7][15] ) );
  LHQD1BWP \vrf/regTable_reg[7][16]  ( .E(n3583), .D(\vrf/N34 ), .Q(
        \vrf/regTable[7][16] ) );
  LHQD1BWP \vrf/regTable_reg[7][17]  ( .E(n3583), .D(\vrf/N35 ), .Q(
        \vrf/regTable[7][17] ) );
  LHQD1BWP \vrf/regTable_reg[7][18]  ( .E(n3583), .D(\vrf/N36 ), .Q(
        \vrf/regTable[7][18] ) );
  LHQD1BWP \vrf/regTable_reg[7][19]  ( .E(n3583), .D(\vrf/N37 ), .Q(
        \vrf/regTable[7][19] ) );
  LHQD1BWP \vrf/regTable_reg[7][20]  ( .E(n3583), .D(\vrf/N38 ), .Q(
        \vrf/regTable[7][20] ) );
  LHQD1BWP \vrf/regTable_reg[7][21]  ( .E(n3583), .D(\vrf/N39 ), .Q(
        \vrf/regTable[7][21] ) );
  LHQD1BWP \vrf/regTable_reg[7][22]  ( .E(n3583), .D(\vrf/N40 ), .Q(
        \vrf/regTable[7][22] ) );
  LHQD1BWP \vrf/regTable_reg[7][23]  ( .E(n3583), .D(\vrf/N41 ), .Q(
        \vrf/regTable[7][23] ) );
  LHQD1BWP \vrf/regTable_reg[7][24]  ( .E(n3583), .D(\vrf/N42 ), .Q(
        \vrf/regTable[7][24] ) );
  LHQD1BWP \vrf/regTable_reg[7][25]  ( .E(n3583), .D(\vrf/N43 ), .Q(
        \vrf/regTable[7][25] ) );
  LHQD1BWP \vrf/regTable_reg[7][26]  ( .E(n3583), .D(\vrf/N44 ), .Q(
        \vrf/regTable[7][26] ) );
  LHQD1BWP \vrf/regTable_reg[7][27]  ( .E(n3583), .D(\vrf/N45 ), .Q(
        \vrf/regTable[7][27] ) );
  LHQD1BWP \vrf/regTable_reg[7][28]  ( .E(n3583), .D(\vrf/N46 ), .Q(
        \vrf/regTable[7][28] ) );
  LHQD1BWP \vrf/regTable_reg[7][29]  ( .E(n3583), .D(\vrf/N47 ), .Q(
        \vrf/regTable[7][29] ) );
  LHQD1BWP \vrf/regTable_reg[7][30]  ( .E(n3583), .D(\vrf/N48 ), .Q(
        \vrf/regTable[7][30] ) );
  LHQD1BWP \vrf/regTable_reg[7][31]  ( .E(n3583), .D(\vrf/N49 ), .Q(
        \vrf/regTable[7][31] ) );
  LHQD1BWP \vrf/regTable_reg[7][32]  ( .E(n3583), .D(\vrf/N50 ), .Q(
        \vrf/regTable[7][32] ) );
  LHQD1BWP \vrf/regTable_reg[7][33]  ( .E(n3583), .D(\vrf/N51 ), .Q(
        \vrf/regTable[7][33] ) );
  LHQD1BWP \vrf/regTable_reg[7][34]  ( .E(n3583), .D(\vrf/N52 ), .Q(
        \vrf/regTable[7][34] ) );
  LHQD1BWP \vrf/regTable_reg[7][35]  ( .E(n3583), .D(\vrf/N53 ), .Q(
        \vrf/regTable[7][35] ) );
  LHQD1BWP \vrf/regTable_reg[7][36]  ( .E(n3583), .D(\vrf/N54 ), .Q(
        \vrf/regTable[7][36] ) );
  LHQD1BWP \vrf/regTable_reg[7][37]  ( .E(n3583), .D(\vrf/N55 ), .Q(
        \vrf/regTable[7][37] ) );
  LHQD1BWP \vrf/regTable_reg[7][38]  ( .E(n3583), .D(\vrf/N56 ), .Q(
        \vrf/regTable[7][38] ) );
  LHQD1BWP \vrf/regTable_reg[7][39]  ( .E(n3583), .D(\vrf/N57 ), .Q(
        \vrf/regTable[7][39] ) );
  LHQD1BWP \vrf/regTable_reg[7][40]  ( .E(n3583), .D(\vrf/N58 ), .Q(
        \vrf/regTable[7][40] ) );
  LHQD1BWP \vrf/regTable_reg[7][41]  ( .E(n3583), .D(\vrf/N59 ), .Q(
        \vrf/regTable[7][41] ) );
  LHQD1BWP \vrf/regTable_reg[7][42]  ( .E(n3583), .D(\vrf/N60 ), .Q(
        \vrf/regTable[7][42] ) );
  LHQD1BWP \vrf/regTable_reg[7][43]  ( .E(n3583), .D(\vrf/N61 ), .Q(
        \vrf/regTable[7][43] ) );
  LHQD1BWP \vrf/regTable_reg[7][44]  ( .E(n3583), .D(\vrf/N62 ), .Q(
        \vrf/regTable[7][44] ) );
  LHQD1BWP \vrf/regTable_reg[7][45]  ( .E(n3583), .D(\vrf/N63 ), .Q(
        \vrf/regTable[7][45] ) );
  LHQD1BWP \vrf/regTable_reg[7][46]  ( .E(n3583), .D(\vrf/N64 ), .Q(
        \vrf/regTable[7][46] ) );
  LHQD1BWP \vrf/regTable_reg[7][47]  ( .E(n3583), .D(\vrf/N65 ), .Q(
        \vrf/regTable[7][47] ) );
  LHQD1BWP \vrf/regTable_reg[7][48]  ( .E(n3583), .D(\vrf/N66 ), .Q(
        \vrf/regTable[7][48] ) );
  LHQD1BWP \vrf/regTable_reg[7][49]  ( .E(n3583), .D(\vrf/N67 ), .Q(
        \vrf/regTable[7][49] ) );
  LHQD1BWP \vrf/regTable_reg[7][50]  ( .E(n3583), .D(\vrf/N68 ), .Q(
        \vrf/regTable[7][50] ) );
  LHQD1BWP \vrf/regTable_reg[7][51]  ( .E(n3583), .D(\vrf/N69 ), .Q(
        \vrf/regTable[7][51] ) );
  LHQD1BWP \vrf/regTable_reg[7][52]  ( .E(n3583), .D(\vrf/N70 ), .Q(
        \vrf/regTable[7][52] ) );
  LHQD1BWP \vrf/regTable_reg[7][53]  ( .E(n3583), .D(\vrf/N71 ), .Q(
        \vrf/regTable[7][53] ) );
  LHQD1BWP \vrf/regTable_reg[7][54]  ( .E(n3583), .D(\vrf/N72 ), .Q(
        \vrf/regTable[7][54] ) );
  LHQD1BWP \vrf/regTable_reg[7][55]  ( .E(n3583), .D(\vrf/N73 ), .Q(
        \vrf/regTable[7][55] ) );
  LHQD1BWP \vrf/regTable_reg[7][56]  ( .E(n3583), .D(\vrf/N74 ), .Q(
        \vrf/regTable[7][56] ) );
  LHQD1BWP \vrf/regTable_reg[7][57]  ( .E(n3583), .D(\vrf/N75 ), .Q(
        \vrf/regTable[7][57] ) );
  LHQD1BWP \vrf/regTable_reg[7][58]  ( .E(n3583), .D(\vrf/N76 ), .Q(
        \vrf/regTable[7][58] ) );
  LHQD1BWP \vrf/regTable_reg[7][59]  ( .E(n3583), .D(\vrf/N77 ), .Q(
        \vrf/regTable[7][59] ) );
  LHQD1BWP \vrf/regTable_reg[7][60]  ( .E(n3583), .D(\vrf/N78 ), .Q(
        \vrf/regTable[7][60] ) );
  LHQD1BWP \vrf/regTable_reg[7][61]  ( .E(n3583), .D(\vrf/N79 ), .Q(
        \vrf/regTable[7][61] ) );
  LHQD1BWP \vrf/regTable_reg[7][62]  ( .E(n3583), .D(\vrf/N80 ), .Q(
        \vrf/regTable[7][62] ) );
  LHQD1BWP \vrf/regTable_reg[7][63]  ( .E(n3583), .D(\vrf/N81 ), .Q(
        \vrf/regTable[7][63] ) );
  LHQD1BWP \vrf/regTable_reg[7][64]  ( .E(n3583), .D(\vrf/N82 ), .Q(
        \vrf/regTable[7][64] ) );
  LHQD1BWP \vrf/regTable_reg[7][65]  ( .E(n3583), .D(\vrf/N83 ), .Q(
        \vrf/regTable[7][65] ) );
  LHQD1BWP \vrf/regTable_reg[7][66]  ( .E(n3583), .D(\vrf/N84 ), .Q(
        \vrf/regTable[7][66] ) );
  LHQD1BWP \vrf/regTable_reg[7][67]  ( .E(n3583), .D(\vrf/N85 ), .Q(
        \vrf/regTable[7][67] ) );
  LHQD1BWP \vrf/regTable_reg[7][68]  ( .E(n3583), .D(\vrf/N86 ), .Q(
        \vrf/regTable[7][68] ) );
  LHQD1BWP \vrf/regTable_reg[7][69]  ( .E(n3583), .D(\vrf/N87 ), .Q(
        \vrf/regTable[7][69] ) );
  LHQD1BWP \vrf/regTable_reg[7][70]  ( .E(n3583), .D(\vrf/N88 ), .Q(
        \vrf/regTable[7][70] ) );
  LHQD1BWP \vrf/regTable_reg[7][71]  ( .E(n3583), .D(\vrf/N89 ), .Q(
        \vrf/regTable[7][71] ) );
  LHQD1BWP \vrf/regTable_reg[7][72]  ( .E(n3583), .D(\vrf/N90 ), .Q(
        \vrf/regTable[7][72] ) );
  LHQD1BWP \vrf/regTable_reg[7][73]  ( .E(n3583), .D(\vrf/N91 ), .Q(
        \vrf/regTable[7][73] ) );
  LHQD1BWP \vrf/regTable_reg[7][74]  ( .E(n3583), .D(\vrf/N92 ), .Q(
        \vrf/regTable[7][74] ) );
  LHQD1BWP \vrf/regTable_reg[7][75]  ( .E(n3583), .D(\vrf/N93 ), .Q(
        \vrf/regTable[7][75] ) );
  LHQD1BWP \vrf/regTable_reg[7][76]  ( .E(n3583), .D(\vrf/N94 ), .Q(
        \vrf/regTable[7][76] ) );
  LHQD1BWP \vrf/regTable_reg[7][77]  ( .E(n3583), .D(\vrf/N95 ), .Q(
        \vrf/regTable[7][77] ) );
  LHQD1BWP \vrf/regTable_reg[7][78]  ( .E(n3583), .D(\vrf/N96 ), .Q(
        \vrf/regTable[7][78] ) );
  LHQD1BWP \vrf/regTable_reg[7][79]  ( .E(n3583), .D(\vrf/N97 ), .Q(
        \vrf/regTable[7][79] ) );
  LHQD1BWP \vrf/regTable_reg[7][80]  ( .E(n3583), .D(\vrf/N98 ), .Q(
        \vrf/regTable[7][80] ) );
  LHQD1BWP \vrf/regTable_reg[7][81]  ( .E(n3583), .D(\vrf/N99 ), .Q(
        \vrf/regTable[7][81] ) );
  LHQD1BWP \vrf/regTable_reg[7][82]  ( .E(n3583), .D(\vrf/N100 ), .Q(
        \vrf/regTable[7][82] ) );
  LHQD1BWP \vrf/regTable_reg[7][83]  ( .E(n3583), .D(\vrf/N101 ), .Q(
        \vrf/regTable[7][83] ) );
  LHQD1BWP \vrf/regTable_reg[7][84]  ( .E(n3583), .D(\vrf/N102 ), .Q(
        \vrf/regTable[7][84] ) );
  LHQD1BWP \vrf/regTable_reg[7][85]  ( .E(n3583), .D(\vrf/N103 ), .Q(
        \vrf/regTable[7][85] ) );
  LHQD1BWP \vrf/regTable_reg[7][86]  ( .E(n3583), .D(\vrf/N104 ), .Q(
        \vrf/regTable[7][86] ) );
  LHQD1BWP \vrf/regTable_reg[7][87]  ( .E(n3583), .D(\vrf/N105 ), .Q(
        \vrf/regTable[7][87] ) );
  LHQD1BWP \vrf/regTable_reg[7][88]  ( .E(n3583), .D(\vrf/N106 ), .Q(
        \vrf/regTable[7][88] ) );
  LHQD1BWP \vrf/regTable_reg[7][89]  ( .E(n3583), .D(\vrf/N107 ), .Q(
        \vrf/regTable[7][89] ) );
  LHQD1BWP \vrf/regTable_reg[7][90]  ( .E(n3583), .D(\vrf/N108 ), .Q(
        \vrf/regTable[7][90] ) );
  LHQD1BWP \vrf/regTable_reg[7][91]  ( .E(n3583), .D(\vrf/N109 ), .Q(
        \vrf/regTable[7][91] ) );
  LHQD1BWP \vrf/regTable_reg[7][92]  ( .E(n3583), .D(\vrf/N110 ), .Q(
        \vrf/regTable[7][92] ) );
  LHQD1BWP \vrf/regTable_reg[7][93]  ( .E(n3583), .D(\vrf/N111 ), .Q(
        \vrf/regTable[7][93] ) );
  LHQD1BWP \vrf/regTable_reg[7][94]  ( .E(n3583), .D(\vrf/N112 ), .Q(
        \vrf/regTable[7][94] ) );
  LHQD1BWP \vrf/regTable_reg[7][95]  ( .E(n3583), .D(\vrf/N113 ), .Q(
        \vrf/regTable[7][95] ) );
  LHQD1BWP \vrf/regTable_reg[7][96]  ( .E(n3583), .D(\vrf/N114 ), .Q(
        \vrf/regTable[7][96] ) );
  LHQD1BWP \vrf/regTable_reg[7][97]  ( .E(n3583), .D(\vrf/N115 ), .Q(
        \vrf/regTable[7][97] ) );
  LHQD1BWP \vrf/regTable_reg[7][98]  ( .E(n3583), .D(\vrf/N116 ), .Q(
        \vrf/regTable[7][98] ) );
  LHQD1BWP \vrf/regTable_reg[7][99]  ( .E(n3583), .D(\vrf/N118 ), .Q(
        \vrf/regTable[7][99] ) );
  LHQD1BWP \vrf/regTable_reg[7][100]  ( .E(n3583), .D(\vrf/N119 ), .Q(
        \vrf/regTable[7][100] ) );
  LHQD1BWP \vrf/regTable_reg[7][101]  ( .E(n3583), .D(\vrf/N120 ), .Q(
        \vrf/regTable[7][101] ) );
  LHQD1BWP \vrf/regTable_reg[7][102]  ( .E(n3583), .D(\vrf/N121 ), .Q(
        \vrf/regTable[7][102] ) );
  LHQD1BWP \vrf/regTable_reg[7][103]  ( .E(n3583), .D(\vrf/N122 ), .Q(
        \vrf/regTable[7][103] ) );
  LHQD1BWP \vrf/regTable_reg[7][104]  ( .E(n3583), .D(\vrf/N123 ), .Q(
        \vrf/regTable[7][104] ) );
  LHQD1BWP \vrf/regTable_reg[7][105]  ( .E(n3583), .D(\vrf/N124 ), .Q(
        \vrf/regTable[7][105] ) );
  LHQD1BWP \vrf/regTable_reg[7][106]  ( .E(n3583), .D(\vrf/N125 ), .Q(
        \vrf/regTable[7][106] ) );
  LHQD1BWP \vrf/regTable_reg[7][107]  ( .E(n3583), .D(\vrf/N126 ), .Q(
        \vrf/regTable[7][107] ) );
  LHQD1BWP \vrf/regTable_reg[7][108]  ( .E(n3583), .D(\vrf/N127 ), .Q(
        \vrf/regTable[7][108] ) );
  LHQD1BWP \vrf/regTable_reg[7][109]  ( .E(n3583), .D(\vrf/N128 ), .Q(
        \vrf/regTable[7][109] ) );
  LHQD1BWP \vrf/regTable_reg[7][110]  ( .E(n3583), .D(\vrf/N129 ), .Q(
        \vrf/regTable[7][110] ) );
  LHQD1BWP \vrf/regTable_reg[7][111]  ( .E(n3583), .D(\vrf/N130 ), .Q(
        \vrf/regTable[7][111] ) );
  LHQD1BWP \vrf/regTable_reg[7][112]  ( .E(n3583), .D(\vrf/N131 ), .Q(
        \vrf/regTable[7][112] ) );
  LHQD1BWP \vrf/regTable_reg[7][113]  ( .E(n3583), .D(\vrf/N132 ), .Q(
        \vrf/regTable[7][113] ) );
  LHQD1BWP \vrf/regTable_reg[7][114]  ( .E(n3583), .D(\vrf/N133 ), .Q(
        \vrf/regTable[7][114] ) );
  LHQD1BWP \vrf/regTable_reg[7][115]  ( .E(n3583), .D(\vrf/N134 ), .Q(
        \vrf/regTable[7][115] ) );
  LHQD1BWP \vrf/regTable_reg[7][116]  ( .E(n3583), .D(\vrf/N135 ), .Q(
        \vrf/regTable[7][116] ) );
  LHQD1BWP \vrf/regTable_reg[7][117]  ( .E(n3583), .D(\vrf/N136 ), .Q(
        \vrf/regTable[7][117] ) );
  LHQD1BWP \vrf/regTable_reg[7][118]  ( .E(n3583), .D(\vrf/N137 ), .Q(
        \vrf/regTable[7][118] ) );
  LHQD1BWP \vrf/regTable_reg[7][119]  ( .E(n3583), .D(\vrf/N138 ), .Q(
        \vrf/regTable[7][119] ) );
  LHQD1BWP \vrf/regTable_reg[7][120]  ( .E(n3583), .D(\vrf/N139 ), .Q(
        \vrf/regTable[7][120] ) );
  LHQD1BWP \vrf/regTable_reg[7][121]  ( .E(n3583), .D(\vrf/N140 ), .Q(
        \vrf/regTable[7][121] ) );
  LHQD1BWP \vrf/regTable_reg[7][122]  ( .E(n3583), .D(\vrf/N141 ), .Q(
        \vrf/regTable[7][122] ) );
  LHQD1BWP \vrf/regTable_reg[7][123]  ( .E(n3583), .D(\vrf/N142 ), .Q(
        \vrf/regTable[7][123] ) );
  LHQD1BWP \vrf/regTable_reg[7][124]  ( .E(n3583), .D(\vrf/N143 ), .Q(
        \vrf/regTable[7][124] ) );
  LHQD1BWP \vrf/regTable_reg[7][125]  ( .E(n3583), .D(\vrf/N144 ), .Q(
        \vrf/regTable[7][125] ) );
  LHQD1BWP \vrf/regTable_reg[7][126]  ( .E(n3583), .D(\vrf/N145 ), .Q(
        \vrf/regTable[7][126] ) );
  LHQD1BWP \vrf/regTable_reg[7][127]  ( .E(n3583), .D(\vrf/N146 ), .Q(
        \vrf/regTable[7][127] ) );
  LHQD1BWP \vrf/regTable_reg[7][128]  ( .E(n3583), .D(\vrf/N147 ), .Q(
        \vrf/regTable[7][128] ) );
  LHQD1BWP \vrf/regTable_reg[7][129]  ( .E(n3583), .D(\vrf/N148 ), .Q(
        \vrf/regTable[7][129] ) );
  LHQD1BWP \vrf/regTable_reg[7][130]  ( .E(n3583), .D(\vrf/N149 ), .Q(
        \vrf/regTable[7][130] ) );
  LHQD1BWP \vrf/regTable_reg[7][131]  ( .E(n3583), .D(\vrf/N150 ), .Q(
        \vrf/regTable[7][131] ) );
  LHQD1BWP \vrf/regTable_reg[7][132]  ( .E(n3583), .D(\vrf/N151 ), .Q(
        \vrf/regTable[7][132] ) );
  LHQD1BWP \vrf/regTable_reg[7][133]  ( .E(n3583), .D(\vrf/N152 ), .Q(
        \vrf/regTable[7][133] ) );
  LHQD1BWP \vrf/regTable_reg[7][134]  ( .E(n3583), .D(\vrf/N153 ), .Q(
        \vrf/regTable[7][134] ) );
  LHQD1BWP \vrf/regTable_reg[7][135]  ( .E(n3583), .D(\vrf/N154 ), .Q(
        \vrf/regTable[7][135] ) );
  LHQD1BWP \vrf/regTable_reg[7][136]  ( .E(n3583), .D(\vrf/N155 ), .Q(
        \vrf/regTable[7][136] ) );
  LHQD1BWP \vrf/regTable_reg[7][137]  ( .E(\vrf/N217 ), .D(\vrf/N156 ), .Q(
        \vrf/regTable[7][137] ) );
  LHQD1BWP \vrf/regTable_reg[7][138]  ( .E(n3583), .D(\vrf/N157 ), .Q(
        \vrf/regTable[7][138] ) );
  LHQD1BWP \vrf/regTable_reg[7][139]  ( .E(\vrf/N217 ), .D(\vrf/N158 ), .Q(
        \vrf/regTable[7][139] ) );
  LHQD1BWP \vrf/regTable_reg[7][140]  ( .E(n3583), .D(\vrf/N159 ), .Q(
        \vrf/regTable[7][140] ) );
  LHQD1BWP \vrf/regTable_reg[7][141]  ( .E(\vrf/N217 ), .D(\vrf/N160 ), .Q(
        \vrf/regTable[7][141] ) );
  LHQD1BWP \vrf/regTable_reg[7][142]  ( .E(n3583), .D(\vrf/N161 ), .Q(
        \vrf/regTable[7][142] ) );
  LHQD1BWP \vrf/regTable_reg[7][143]  ( .E(\vrf/N217 ), .D(\vrf/N162 ), .Q(
        \vrf/regTable[7][143] ) );
  LHQD1BWP \vrf/regTable_reg[7][144]  ( .E(n3583), .D(\vrf/N163 ), .Q(
        \vrf/regTable[7][144] ) );
  LHQD1BWP \vrf/regTable_reg[7][145]  ( .E(\vrf/N217 ), .D(\vrf/N164 ), .Q(
        \vrf/regTable[7][145] ) );
  LHQD1BWP \vrf/regTable_reg[7][146]  ( .E(n3583), .D(\vrf/N165 ), .Q(
        \vrf/regTable[7][146] ) );
  LHQD1BWP \vrf/regTable_reg[7][147]  ( .E(\vrf/N217 ), .D(\vrf/N166 ), .Q(
        \vrf/regTable[7][147] ) );
  LHQD1BWP \vrf/regTable_reg[7][148]  ( .E(n3583), .D(\vrf/N167 ), .Q(
        \vrf/regTable[7][148] ) );
  LHQD1BWP \vrf/regTable_reg[7][149]  ( .E(n3583), .D(\vrf/N168 ), .Q(
        \vrf/regTable[7][149] ) );
  LHQD1BWP \vrf/regTable_reg[7][150]  ( .E(n3583), .D(\vrf/N169 ), .Q(
        \vrf/regTable[7][150] ) );
  LHQD1BWP \vrf/regTable_reg[7][151]  ( .E(\vrf/N217 ), .D(\vrf/N170 ), .Q(
        \vrf/regTable[7][151] ) );
  LHQD1BWP \vrf/regTable_reg[7][152]  ( .E(n3583), .D(\vrf/N171 ), .Q(
        \vrf/regTable[7][152] ) );
  LHQD1BWP \vrf/regTable_reg[7][153]  ( .E(n3583), .D(\vrf/N172 ), .Q(
        \vrf/regTable[7][153] ) );
  LHQD1BWP \vrf/regTable_reg[7][154]  ( .E(n3583), .D(\vrf/N173 ), .Q(
        \vrf/regTable[7][154] ) );
  LHQD1BWP \vrf/regTable_reg[7][155]  ( .E(\vrf/N217 ), .D(\vrf/N174 ), .Q(
        \vrf/regTable[7][155] ) );
  LHQD1BWP \vrf/regTable_reg[7][156]  ( .E(n3583), .D(\vrf/N175 ), .Q(
        \vrf/regTable[7][156] ) );
  LHQD1BWP \vrf/regTable_reg[7][157]  ( .E(n3583), .D(\vrf/N176 ), .Q(
        \vrf/regTable[7][157] ) );
  LHQD1BWP \vrf/regTable_reg[7][158]  ( .E(n3583), .D(\vrf/N177 ), .Q(
        \vrf/regTable[7][158] ) );
  LHQD1BWP \vrf/regTable_reg[7][159]  ( .E(n3583), .D(\vrf/N178 ), .Q(
        \vrf/regTable[7][159] ) );
  LHQD1BWP \vrf/regTable_reg[7][160]  ( .E(\vrf/N217 ), .D(\vrf/N179 ), .Q(
        \vrf/regTable[7][160] ) );
  LHQD1BWP \vrf/regTable_reg[7][161]  ( .E(n3583), .D(\vrf/N180 ), .Q(
        \vrf/regTable[7][161] ) );
  LHQD1BWP \vrf/regTable_reg[7][162]  ( .E(n3583), .D(\vrf/N181 ), .Q(
        \vrf/regTable[7][162] ) );
  LHQD1BWP \vrf/regTable_reg[7][163]  ( .E(n3583), .D(\vrf/N182 ), .Q(
        \vrf/regTable[7][163] ) );
  LHQD1BWP \vrf/regTable_reg[7][164]  ( .E(\vrf/N217 ), .D(\vrf/N183 ), .Q(
        \vrf/regTable[7][164] ) );
  LHQD1BWP \vrf/regTable_reg[7][165]  ( .E(n3583), .D(\vrf/N184 ), .Q(
        \vrf/regTable[7][165] ) );
  LHQD1BWP \vrf/regTable_reg[7][166]  ( .E(n3583), .D(\vrf/N185 ), .Q(
        \vrf/regTable[7][166] ) );
  LHQD1BWP \vrf/regTable_reg[7][167]  ( .E(n3583), .D(\vrf/N186 ), .Q(
        \vrf/regTable[7][167] ) );
  LHQD1BWP \vrf/regTable_reg[7][168]  ( .E(\vrf/N217 ), .D(\vrf/N187 ), .Q(
        \vrf/regTable[7][168] ) );
  LHQD1BWP \vrf/regTable_reg[7][169]  ( .E(n3583), .D(\vrf/N188 ), .Q(
        \vrf/regTable[7][169] ) );
  LHQD1BWP \vrf/regTable_reg[7][170]  ( .E(n3583), .D(\vrf/N189 ), .Q(
        \vrf/regTable[7][170] ) );
  LHQD1BWP \vrf/regTable_reg[7][171]  ( .E(n3583), .D(\vrf/N190 ), .Q(
        \vrf/regTable[7][171] ) );
  LHQD1BWP \vrf/regTable_reg[7][172]  ( .E(n3583), .D(\vrf/N191 ), .Q(
        \vrf/regTable[7][172] ) );
  LHQD1BWP \vrf/regTable_reg[7][173]  ( .E(n3583), .D(\vrf/N192 ), .Q(
        \vrf/regTable[7][173] ) );
  LHQD1BWP \vrf/regTable_reg[7][174]  ( .E(\vrf/N217 ), .D(\vrf/N193 ), .Q(
        \vrf/regTable[7][174] ) );
  LHQD1BWP \vrf/regTable_reg[7][175]  ( .E(n3583), .D(\vrf/N194 ), .Q(
        \vrf/regTable[7][175] ) );
  LHQD1BWP \vrf/regTable_reg[7][176]  ( .E(n3583), .D(\vrf/N195 ), .Q(
        \vrf/regTable[7][176] ) );
  LHQD1BWP \vrf/regTable_reg[7][177]  ( .E(n3583), .D(\vrf/N196 ), .Q(
        \vrf/regTable[7][177] ) );
  LHQD1BWP \vrf/regTable_reg[7][178]  ( .E(n3583), .D(\vrf/N197 ), .Q(
        \vrf/regTable[7][178] ) );
  LHQD1BWP \vrf/regTable_reg[7][179]  ( .E(\vrf/N217 ), .D(\vrf/N198 ), .Q(
        \vrf/regTable[7][179] ) );
  LHQD1BWP \vrf/regTable_reg[7][180]  ( .E(n3583), .D(\vrf/N199 ), .Q(
        \vrf/regTable[7][180] ) );
  LHQD1BWP \vrf/regTable_reg[7][181]  ( .E(n3583), .D(\vrf/N200 ), .Q(
        \vrf/regTable[7][181] ) );
  LHQD1BWP \vrf/regTable_reg[7][182]  ( .E(n3583), .D(\vrf/N201 ), .Q(
        \vrf/regTable[7][182] ) );
  LHQD1BWP \vrf/regTable_reg[7][183]  ( .E(n3583), .D(\vrf/N202 ), .Q(
        \vrf/regTable[7][183] ) );
  LHQD1BWP \vrf/regTable_reg[7][184]  ( .E(n3583), .D(\vrf/N203 ), .Q(
        \vrf/regTable[7][184] ) );
  LHQD1BWP \vrf/regTable_reg[7][185]  ( .E(n3583), .D(\vrf/N204 ), .Q(
        \vrf/regTable[7][185] ) );
  LHQD1BWP \vrf/regTable_reg[7][186]  ( .E(n3583), .D(\vrf/N205 ), .Q(
        \vrf/regTable[7][186] ) );
  LHQD1BWP \vrf/regTable_reg[7][187]  ( .E(n3583), .D(\vrf/N206 ), .Q(
        \vrf/regTable[7][187] ) );
  LHQD1BWP \vrf/regTable_reg[7][188]  ( .E(n3583), .D(\vrf/N207 ), .Q(
        \vrf/regTable[7][188] ) );
  LHQD1BWP \vrf/regTable_reg[7][189]  ( .E(\vrf/N217 ), .D(\vrf/N208 ), .Q(
        \vrf/regTable[7][189] ) );
  LHQD1BWP \vrf/regTable_reg[7][190]  ( .E(n3583), .D(\vrf/N209 ), .Q(
        \vrf/regTable[7][190] ) );
  LHQD1BWP \vrf/regTable_reg[7][191]  ( .E(n3583), .D(\vrf/N210 ), .Q(
        \vrf/regTable[7][191] ) );
  LHQD1BWP \vrf/regTable_reg[7][192]  ( .E(n3583), .D(\vrf/N211 ), .Q(
        \vrf/regTable[7][192] ) );
  LHQD1BWP \vrf/regTable_reg[7][193]  ( .E(n3583), .D(\vrf/N212 ), .Q(
        \vrf/regTable[7][193] ) );
  LHQD1BWP \vrf/regTable_reg[7][194]  ( .E(\vrf/N217 ), .D(\vrf/N213 ), .Q(
        \vrf/regTable[7][194] ) );
  LHQD1BWP \vrf/regTable_reg[7][195]  ( .E(\vrf/N217 ), .D(\vrf/N214 ), .Q(
        \vrf/regTable[7][195] ) );
  LHQD1BWP \vrf/regTable_reg[7][196]  ( .E(n3583), .D(\vrf/N215 ), .Q(
        \vrf/regTable[7][196] ) );
  LHQD1BWP \vrf/regTable_reg[7][197]  ( .E(n3583), .D(\vrf/N216 ), .Q(
        \vrf/regTable[7][197] ) );
  LHQD1BWP \vrf/regTable_reg[7][198]  ( .E(n3583), .D(\vrf/N218 ), .Q(
        \vrf/regTable[7][198] ) );
  LHQD1BWP \vrf/regTable_reg[7][199]  ( .E(n3583), .D(\vrf/N219 ), .Q(
        \vrf/regTable[7][199] ) );
  LHQD1BWP \vrf/regTable_reg[7][200]  ( .E(n3583), .D(\vrf/N220 ), .Q(
        \vrf/regTable[7][200] ) );
  LHQD1BWP \vrf/regTable_reg[7][201]  ( .E(\vrf/N217 ), .D(\vrf/N221 ), .Q(
        \vrf/regTable[7][201] ) );
  LHQD1BWP \vrf/regTable_reg[7][202]  ( .E(n3583), .D(\vrf/N222 ), .Q(
        \vrf/regTable[7][202] ) );
  LHQD1BWP \vrf/regTable_reg[7][203]  ( .E(n3583), .D(\vrf/N223 ), .Q(
        \vrf/regTable[7][203] ) );
  LHQD1BWP \vrf/regTable_reg[7][204]  ( .E(\vrf/N217 ), .D(\vrf/N224 ), .Q(
        \vrf/regTable[7][204] ) );
  LHQD1BWP \vrf/regTable_reg[7][205]  ( .E(n3583), .D(\vrf/N225 ), .Q(
        \vrf/regTable[7][205] ) );
  LHQD1BWP \vrf/regTable_reg[7][206]  ( .E(\vrf/N217 ), .D(\vrf/N226 ), .Q(
        \vrf/regTable[7][206] ) );
  LHQD1BWP \vrf/regTable_reg[7][207]  ( .E(n3583), .D(\vrf/N227 ), .Q(
        \vrf/regTable[7][207] ) );
  LHQD1BWP \vrf/regTable_reg[7][208]  ( .E(n3583), .D(\vrf/N228 ), .Q(
        \vrf/regTable[7][208] ) );
  LHQD1BWP \vrf/regTable_reg[7][209]  ( .E(n3583), .D(\vrf/N229 ), .Q(
        \vrf/regTable[7][209] ) );
  LHQD1BWP \vrf/regTable_reg[7][210]  ( .E(n3583), .D(\vrf/N230 ), .Q(
        \vrf/regTable[7][210] ) );
  LHQD1BWP \vrf/regTable_reg[7][211]  ( .E(n3583), .D(\vrf/N231 ), .Q(
        \vrf/regTable[7][211] ) );
  LHQD1BWP \vrf/regTable_reg[7][212]  ( .E(n3583), .D(\vrf/N232 ), .Q(
        \vrf/regTable[7][212] ) );
  LHQD1BWP \vrf/regTable_reg[7][213]  ( .E(n3583), .D(\vrf/N233 ), .Q(
        \vrf/regTable[7][213] ) );
  LHQD1BWP \vrf/regTable_reg[7][214]  ( .E(n3583), .D(\vrf/N234 ), .Q(
        \vrf/regTable[7][214] ) );
  LHQD1BWP \vrf/regTable_reg[7][215]  ( .E(n3583), .D(\vrf/N235 ), .Q(
        \vrf/regTable[7][215] ) );
  LHQD1BWP \vrf/regTable_reg[7][216]  ( .E(n3583), .D(\vrf/N236 ), .Q(
        \vrf/regTable[7][216] ) );
  LHQD1BWP \vrf/regTable_reg[7][217]  ( .E(n3583), .D(\vrf/N237 ), .Q(
        \vrf/regTable[7][217] ) );
  LHQD1BWP \vrf/regTable_reg[7][218]  ( .E(n3583), .D(\vrf/N238 ), .Q(
        \vrf/regTable[7][218] ) );
  LHQD1BWP \vrf/regTable_reg[7][219]  ( .E(n3583), .D(\vrf/N239 ), .Q(
        \vrf/regTable[7][219] ) );
  LHQD1BWP \vrf/regTable_reg[7][220]  ( .E(n3583), .D(\vrf/N240 ), .Q(
        \vrf/regTable[7][220] ) );
  LHQD1BWP \vrf/regTable_reg[7][221]  ( .E(n3583), .D(\vrf/N241 ), .Q(
        \vrf/regTable[7][221] ) );
  LHQD1BWP \vrf/regTable_reg[7][222]  ( .E(n3583), .D(\vrf/N242 ), .Q(
        \vrf/regTable[7][222] ) );
  LHQD1BWP \vrf/regTable_reg[7][223]  ( .E(\vrf/N217 ), .D(\vrf/N243 ), .Q(
        \vrf/regTable[7][223] ) );
  LHQD1BWP \vrf/regTable_reg[7][224]  ( .E(n3583), .D(\vrf/N244 ), .Q(
        \vrf/regTable[7][224] ) );
  LHQD1BWP \vrf/regTable_reg[7][225]  ( .E(n3583), .D(\vrf/N245 ), .Q(
        \vrf/regTable[7][225] ) );
  LHQD1BWP \vrf/regTable_reg[7][226]  ( .E(n3583), .D(\vrf/N246 ), .Q(
        \vrf/regTable[7][226] ) );
  LHQD1BWP \vrf/regTable_reg[7][227]  ( .E(\vrf/N217 ), .D(\vrf/N247 ), .Q(
        \vrf/regTable[7][227] ) );
  LHQD1BWP \vrf/regTable_reg[7][228]  ( .E(n3583), .D(\vrf/N248 ), .Q(
        \vrf/regTable[7][228] ) );
  LHQD1BWP \vrf/regTable_reg[7][229]  ( .E(n3583), .D(\vrf/N249 ), .Q(
        \vrf/regTable[7][229] ) );
  LHQD1BWP \vrf/regTable_reg[7][230]  ( .E(n3583), .D(\vrf/N250 ), .Q(
        \vrf/regTable[7][230] ) );
  LHQD1BWP \vrf/regTable_reg[7][231]  ( .E(\vrf/N217 ), .D(\vrf/N251 ), .Q(
        \vrf/regTable[7][231] ) );
  LHQD1BWP \vrf/regTable_reg[7][232]  ( .E(n3583), .D(\vrf/N252 ), .Q(
        \vrf/regTable[7][232] ) );
  LHQD1BWP \vrf/regTable_reg[7][233]  ( .E(n3583), .D(\vrf/N253 ), .Q(
        \vrf/regTable[7][233] ) );
  LHQD1BWP \vrf/regTable_reg[7][234]  ( .E(n3583), .D(\vrf/N254 ), .Q(
        \vrf/regTable[7][234] ) );
  LHQD1BWP \vrf/regTable_reg[7][235]  ( .E(n3583), .D(\vrf/N255 ), .Q(
        \vrf/regTable[7][235] ) );
  LHQD1BWP \vrf/regTable_reg[7][236]  ( .E(n3583), .D(\vrf/N256 ), .Q(
        \vrf/regTable[7][236] ) );
  LHQD1BWP \vrf/regTable_reg[7][237]  ( .E(n3583), .D(\vrf/N257 ), .Q(
        \vrf/regTable[7][237] ) );
  LHQD1BWP \vrf/regTable_reg[7][238]  ( .E(n3583), .D(\vrf/N258 ), .Q(
        \vrf/regTable[7][238] ) );
  LHQD1BWP \vrf/regTable_reg[7][239]  ( .E(n3583), .D(\vrf/N259 ), .Q(
        \vrf/regTable[7][239] ) );
  LHQD1BWP \vrf/regTable_reg[7][240]  ( .E(n3583), .D(\vrf/N260 ), .Q(
        \vrf/regTable[7][240] ) );
  LHQD1BWP \vrf/regTable_reg[7][241]  ( .E(n3583), .D(\vrf/N261 ), .Q(
        \vrf/regTable[7][241] ) );
  LHQD1BWP \vrf/regTable_reg[7][242]  ( .E(n3583), .D(\vrf/N262 ), .Q(
        \vrf/regTable[7][242] ) );
  LHQD1BWP \vrf/regTable_reg[7][243]  ( .E(n3583), .D(\vrf/N263 ), .Q(
        \vrf/regTable[7][243] ) );
  LHQD1BWP \vrf/regTable_reg[7][244]  ( .E(n3583), .D(\vrf/N264 ), .Q(
        \vrf/regTable[7][244] ) );
  LHQD1BWP \vrf/regTable_reg[7][245]  ( .E(n3583), .D(\vrf/N265 ), .Q(
        \vrf/regTable[7][245] ) );
  LHQD1BWP \vrf/regTable_reg[7][246]  ( .E(n3583), .D(\vrf/N266 ), .Q(
        \vrf/regTable[7][246] ) );
  LHQD1BWP \vrf/regTable_reg[7][247]  ( .E(n3583), .D(\vrf/N267 ), .Q(
        \vrf/regTable[7][247] ) );
  LHQD1BWP \vrf/regTable_reg[7][248]  ( .E(n3583), .D(\vrf/N268 ), .Q(
        \vrf/regTable[7][248] ) );
  LHQD1BWP \vrf/regTable_reg[7][249]  ( .E(n3583), .D(\vrf/N269 ), .Q(
        \vrf/regTable[7][249] ) );
  LHQD1BWP \vrf/regTable_reg[7][250]  ( .E(n3583), .D(\vrf/N270 ), .Q(
        \vrf/regTable[7][250] ) );
  LHQD1BWP \vrf/regTable_reg[7][251]  ( .E(\vrf/N217 ), .D(\vrf/N271 ), .Q(
        \vrf/regTable[7][251] ) );
  LHQD1BWP \vrf/regTable_reg[7][252]  ( .E(n3583), .D(\vrf/N272 ), .Q(
        \vrf/regTable[7][252] ) );
  LHQD1BWP \vrf/regTable_reg[7][253]  ( .E(n3583), .D(\vrf/N273 ), .Q(
        \vrf/regTable[7][253] ) );
  LHQD1BWP \vrf/regTable_reg[7][254]  ( .E(n3583), .D(\vrf/N274 ), .Q(
        \vrf/regTable[7][254] ) );
  LHQD1BWP \vrf/regTable_reg[7][255]  ( .E(n3583), .D(\vrf/N275 ), .Q(
        \vrf/regTable[7][255] ) );
  LHQD1BWP \vrf/regTable_reg[6][0]  ( .E(n3585), .D(\vrf/N18 ), .Q(
        \vrf/regTable[6][0] ) );
  LHQD1BWP \vrf/regTable_reg[6][1]  ( .E(n3585), .D(\vrf/N19 ), .Q(
        \vrf/regTable[6][1] ) );
  LHQD1BWP \vrf/regTable_reg[6][2]  ( .E(n3585), .D(\vrf/N20 ), .Q(
        \vrf/regTable[6][2] ) );
  LHQD1BWP \vrf/regTable_reg[6][3]  ( .E(n3585), .D(\vrf/N21 ), .Q(
        \vrf/regTable[6][3] ) );
  LHQD1BWP \vrf/regTable_reg[6][4]  ( .E(n3585), .D(\vrf/N22 ), .Q(
        \vrf/regTable[6][4] ) );
  LHQD1BWP \vrf/regTable_reg[6][5]  ( .E(n3585), .D(\vrf/N23 ), .Q(
        \vrf/regTable[6][5] ) );
  LHQD1BWP \vrf/regTable_reg[6][6]  ( .E(n3585), .D(\vrf/N24 ), .Q(
        \vrf/regTable[6][6] ) );
  LHQD1BWP \vrf/regTable_reg[6][7]  ( .E(n3585), .D(\vrf/N25 ), .Q(
        \vrf/regTable[6][7] ) );
  LHQD1BWP \vrf/regTable_reg[6][8]  ( .E(n3585), .D(\vrf/N26 ), .Q(
        \vrf/regTable[6][8] ) );
  LHQD1BWP \vrf/regTable_reg[6][9]  ( .E(n3585), .D(\vrf/N27 ), .Q(
        \vrf/regTable[6][9] ) );
  LHQD1BWP \vrf/regTable_reg[6][10]  ( .E(n3585), .D(\vrf/N28 ), .Q(
        \vrf/regTable[6][10] ) );
  LHQD1BWP \vrf/regTable_reg[6][11]  ( .E(n3585), .D(\vrf/N29 ), .Q(
        \vrf/regTable[6][11] ) );
  LHQD1BWP \vrf/regTable_reg[6][12]  ( .E(n3585), .D(\vrf/N30 ), .Q(
        \vrf/regTable[6][12] ) );
  LHQD1BWP \vrf/regTable_reg[6][13]  ( .E(n3585), .D(\vrf/N31 ), .Q(
        \vrf/regTable[6][13] ) );
  LHQD1BWP \vrf/regTable_reg[6][14]  ( .E(n3585), .D(\vrf/N32 ), .Q(
        \vrf/regTable[6][14] ) );
  LHQD1BWP \vrf/regTable_reg[6][15]  ( .E(n3585), .D(\vrf/N33 ), .Q(
        \vrf/regTable[6][15] ) );
  LHQD1BWP \vrf/regTable_reg[6][16]  ( .E(n3585), .D(\vrf/N34 ), .Q(
        \vrf/regTable[6][16] ) );
  LHQD1BWP \vrf/regTable_reg[6][17]  ( .E(n3585), .D(\vrf/N35 ), .Q(
        \vrf/regTable[6][17] ) );
  LHQD1BWP \vrf/regTable_reg[6][18]  ( .E(n3585), .D(\vrf/N36 ), .Q(
        \vrf/regTable[6][18] ) );
  LHQD1BWP \vrf/regTable_reg[6][19]  ( .E(n3585), .D(\vrf/N37 ), .Q(
        \vrf/regTable[6][19] ) );
  LHQD1BWP \vrf/regTable_reg[6][20]  ( .E(n3585), .D(\vrf/N38 ), .Q(
        \vrf/regTable[6][20] ) );
  LHQD1BWP \vrf/regTable_reg[6][21]  ( .E(n3585), .D(\vrf/N39 ), .Q(
        \vrf/regTable[6][21] ) );
  LHQD1BWP \vrf/regTable_reg[6][22]  ( .E(n3585), .D(\vrf/N40 ), .Q(
        \vrf/regTable[6][22] ) );
  LHQD1BWP \vrf/regTable_reg[6][23]  ( .E(n3585), .D(\vrf/N41 ), .Q(
        \vrf/regTable[6][23] ) );
  LHQD1BWP \vrf/regTable_reg[6][24]  ( .E(n3585), .D(\vrf/N42 ), .Q(
        \vrf/regTable[6][24] ) );
  LHQD1BWP \vrf/regTable_reg[6][25]  ( .E(n3585), .D(\vrf/N43 ), .Q(
        \vrf/regTable[6][25] ) );
  LHQD1BWP \vrf/regTable_reg[6][26]  ( .E(n3585), .D(\vrf/N44 ), .Q(
        \vrf/regTable[6][26] ) );
  LHQD1BWP \vrf/regTable_reg[6][27]  ( .E(n3585), .D(\vrf/N45 ), .Q(
        \vrf/regTable[6][27] ) );
  LHQD1BWP \vrf/regTable_reg[6][28]  ( .E(n3585), .D(\vrf/N46 ), .Q(
        \vrf/regTable[6][28] ) );
  LHQD1BWP \vrf/regTable_reg[6][29]  ( .E(n3585), .D(\vrf/N47 ), .Q(
        \vrf/regTable[6][29] ) );
  LHQD1BWP \vrf/regTable_reg[6][30]  ( .E(n3585), .D(\vrf/N48 ), .Q(
        \vrf/regTable[6][30] ) );
  LHQD1BWP \vrf/regTable_reg[6][31]  ( .E(n3585), .D(\vrf/N49 ), .Q(
        \vrf/regTable[6][31] ) );
  LHQD1BWP \vrf/regTable_reg[6][32]  ( .E(n3585), .D(\vrf/N50 ), .Q(
        \vrf/regTable[6][32] ) );
  LHQD1BWP \vrf/regTable_reg[6][33]  ( .E(n3585), .D(\vrf/N51 ), .Q(
        \vrf/regTable[6][33] ) );
  LHQD1BWP \vrf/regTable_reg[6][34]  ( .E(n3585), .D(\vrf/N52 ), .Q(
        \vrf/regTable[6][34] ) );
  LHQD1BWP \vrf/regTable_reg[6][35]  ( .E(n3585), .D(\vrf/N53 ), .Q(
        \vrf/regTable[6][35] ) );
  LHQD1BWP \vrf/regTable_reg[6][36]  ( .E(n3585), .D(\vrf/N54 ), .Q(
        \vrf/regTable[6][36] ) );
  LHQD1BWP \vrf/regTable_reg[6][37]  ( .E(n3585), .D(\vrf/N55 ), .Q(
        \vrf/regTable[6][37] ) );
  LHQD1BWP \vrf/regTable_reg[6][38]  ( .E(n3585), .D(\vrf/N56 ), .Q(
        \vrf/regTable[6][38] ) );
  LHQD1BWP \vrf/regTable_reg[6][39]  ( .E(n3585), .D(\vrf/N57 ), .Q(
        \vrf/regTable[6][39] ) );
  LHQD1BWP \vrf/regTable_reg[6][40]  ( .E(n3585), .D(\vrf/N58 ), .Q(
        \vrf/regTable[6][40] ) );
  LHQD1BWP \vrf/regTable_reg[6][41]  ( .E(n3585), .D(\vrf/N59 ), .Q(
        \vrf/regTable[6][41] ) );
  LHQD1BWP \vrf/regTable_reg[6][42]  ( .E(n3585), .D(\vrf/N60 ), .Q(
        \vrf/regTable[6][42] ) );
  LHQD1BWP \vrf/regTable_reg[6][43]  ( .E(n3585), .D(\vrf/N61 ), .Q(
        \vrf/regTable[6][43] ) );
  LHQD1BWP \vrf/regTable_reg[6][44]  ( .E(n3585), .D(\vrf/N62 ), .Q(
        \vrf/regTable[6][44] ) );
  LHQD1BWP \vrf/regTable_reg[6][45]  ( .E(n3585), .D(\vrf/N63 ), .Q(
        \vrf/regTable[6][45] ) );
  LHQD1BWP \vrf/regTable_reg[6][46]  ( .E(n3585), .D(\vrf/N64 ), .Q(
        \vrf/regTable[6][46] ) );
  LHQD1BWP \vrf/regTable_reg[6][47]  ( .E(n3585), .D(\vrf/N65 ), .Q(
        \vrf/regTable[6][47] ) );
  LHQD1BWP \vrf/regTable_reg[6][48]  ( .E(n3585), .D(\vrf/N66 ), .Q(
        \vrf/regTable[6][48] ) );
  LHQD1BWP \vrf/regTable_reg[6][49]  ( .E(n3585), .D(\vrf/N67 ), .Q(
        \vrf/regTable[6][49] ) );
  LHQD1BWP \vrf/regTable_reg[6][50]  ( .E(n3585), .D(\vrf/N68 ), .Q(
        \vrf/regTable[6][50] ) );
  LHQD1BWP \vrf/regTable_reg[6][51]  ( .E(n3585), .D(\vrf/N69 ), .Q(
        \vrf/regTable[6][51] ) );
  LHQD1BWP \vrf/regTable_reg[6][52]  ( .E(n3585), .D(\vrf/N70 ), .Q(
        \vrf/regTable[6][52] ) );
  LHQD1BWP \vrf/regTable_reg[6][53]  ( .E(n3585), .D(\vrf/N71 ), .Q(
        \vrf/regTable[6][53] ) );
  LHQD1BWP \vrf/regTable_reg[6][54]  ( .E(n3585), .D(\vrf/N72 ), .Q(
        \vrf/regTable[6][54] ) );
  LHQD1BWP \vrf/regTable_reg[6][55]  ( .E(n3585), .D(\vrf/N73 ), .Q(
        \vrf/regTable[6][55] ) );
  LHQD1BWP \vrf/regTable_reg[6][56]  ( .E(n3585), .D(\vrf/N74 ), .Q(
        \vrf/regTable[6][56] ) );
  LHQD1BWP \vrf/regTable_reg[6][57]  ( .E(n3585), .D(\vrf/N75 ), .Q(
        \vrf/regTable[6][57] ) );
  LHQD1BWP \vrf/regTable_reg[6][58]  ( .E(n3585), .D(\vrf/N76 ), .Q(
        \vrf/regTable[6][58] ) );
  LHQD1BWP \vrf/regTable_reg[6][59]  ( .E(n3585), .D(\vrf/N77 ), .Q(
        \vrf/regTable[6][59] ) );
  LHQD1BWP \vrf/regTable_reg[6][60]  ( .E(n3585), .D(\vrf/N78 ), .Q(
        \vrf/regTable[6][60] ) );
  LHQD1BWP \vrf/regTable_reg[6][61]  ( .E(n3585), .D(\vrf/N79 ), .Q(
        \vrf/regTable[6][61] ) );
  LHQD1BWP \vrf/regTable_reg[6][62]  ( .E(n3585), .D(\vrf/N80 ), .Q(
        \vrf/regTable[6][62] ) );
  LHQD1BWP \vrf/regTable_reg[6][63]  ( .E(n3585), .D(\vrf/N81 ), .Q(
        \vrf/regTable[6][63] ) );
  LHQD1BWP \vrf/regTable_reg[6][64]  ( .E(n3585), .D(\vrf/N82 ), .Q(
        \vrf/regTable[6][64] ) );
  LHQD1BWP \vrf/regTable_reg[6][65]  ( .E(n3585), .D(\vrf/N83 ), .Q(
        \vrf/regTable[6][65] ) );
  LHQD1BWP \vrf/regTable_reg[6][66]  ( .E(n3585), .D(\vrf/N84 ), .Q(
        \vrf/regTable[6][66] ) );
  LHQD1BWP \vrf/regTable_reg[6][67]  ( .E(n3585), .D(\vrf/N85 ), .Q(
        \vrf/regTable[6][67] ) );
  LHQD1BWP \vrf/regTable_reg[6][68]  ( .E(n3585), .D(\vrf/N86 ), .Q(
        \vrf/regTable[6][68] ) );
  LHQD1BWP \vrf/regTable_reg[6][69]  ( .E(n3585), .D(\vrf/N87 ), .Q(
        \vrf/regTable[6][69] ) );
  LHQD1BWP \vrf/regTable_reg[6][70]  ( .E(n3585), .D(\vrf/N88 ), .Q(
        \vrf/regTable[6][70] ) );
  LHQD1BWP \vrf/regTable_reg[6][71]  ( .E(n3585), .D(\vrf/N89 ), .Q(
        \vrf/regTable[6][71] ) );
  LHQD1BWP \vrf/regTable_reg[6][72]  ( .E(n3585), .D(\vrf/N90 ), .Q(
        \vrf/regTable[6][72] ) );
  LHQD1BWP \vrf/regTable_reg[6][73]  ( .E(n3585), .D(\vrf/N91 ), .Q(
        \vrf/regTable[6][73] ) );
  LHQD1BWP \vrf/regTable_reg[6][74]  ( .E(n3585), .D(\vrf/N92 ), .Q(
        \vrf/regTable[6][74] ) );
  LHQD1BWP \vrf/regTable_reg[6][75]  ( .E(n3585), .D(\vrf/N93 ), .Q(
        \vrf/regTable[6][75] ) );
  LHQD1BWP \vrf/regTable_reg[6][76]  ( .E(n3585), .D(\vrf/N94 ), .Q(
        \vrf/regTable[6][76] ) );
  LHQD1BWP \vrf/regTable_reg[6][77]  ( .E(n3585), .D(\vrf/N95 ), .Q(
        \vrf/regTable[6][77] ) );
  LHQD1BWP \vrf/regTable_reg[6][78]  ( .E(n3585), .D(\vrf/N96 ), .Q(
        \vrf/regTable[6][78] ) );
  LHQD1BWP \vrf/regTable_reg[6][79]  ( .E(n3585), .D(\vrf/N97 ), .Q(
        \vrf/regTable[6][79] ) );
  LHQD1BWP \vrf/regTable_reg[6][80]  ( .E(n3585), .D(\vrf/N98 ), .Q(
        \vrf/regTable[6][80] ) );
  LHQD1BWP \vrf/regTable_reg[6][81]  ( .E(n3585), .D(\vrf/N99 ), .Q(
        \vrf/regTable[6][81] ) );
  LHQD1BWP \vrf/regTable_reg[6][82]  ( .E(n3585), .D(\vrf/N100 ), .Q(
        \vrf/regTable[6][82] ) );
  LHQD1BWP \vrf/regTable_reg[6][83]  ( .E(n3585), .D(\vrf/N101 ), .Q(
        \vrf/regTable[6][83] ) );
  LHQD1BWP \vrf/regTable_reg[6][84]  ( .E(n3585), .D(\vrf/N102 ), .Q(
        \vrf/regTable[6][84] ) );
  LHQD1BWP \vrf/regTable_reg[6][85]  ( .E(n3585), .D(\vrf/N103 ), .Q(
        \vrf/regTable[6][85] ) );
  LHQD1BWP \vrf/regTable_reg[6][86]  ( .E(n3585), .D(\vrf/N104 ), .Q(
        \vrf/regTable[6][86] ) );
  LHQD1BWP \vrf/regTable_reg[6][87]  ( .E(n3585), .D(\vrf/N105 ), .Q(
        \vrf/regTable[6][87] ) );
  LHQD1BWP \vrf/regTable_reg[6][88]  ( .E(n3585), .D(\vrf/N106 ), .Q(
        \vrf/regTable[6][88] ) );
  LHQD1BWP \vrf/regTable_reg[6][89]  ( .E(n3585), .D(\vrf/N107 ), .Q(
        \vrf/regTable[6][89] ) );
  LHQD1BWP \vrf/regTable_reg[6][90]  ( .E(n3585), .D(\vrf/N108 ), .Q(
        \vrf/regTable[6][90] ) );
  LHQD1BWP \vrf/regTable_reg[6][91]  ( .E(n3585), .D(\vrf/N109 ), .Q(
        \vrf/regTable[6][91] ) );
  LHQD1BWP \vrf/regTable_reg[6][92]  ( .E(n3585), .D(\vrf/N110 ), .Q(
        \vrf/regTable[6][92] ) );
  LHQD1BWP \vrf/regTable_reg[6][93]  ( .E(n3585), .D(\vrf/N111 ), .Q(
        \vrf/regTable[6][93] ) );
  LHQD1BWP \vrf/regTable_reg[6][94]  ( .E(n3585), .D(\vrf/N112 ), .Q(
        \vrf/regTable[6][94] ) );
  LHQD1BWP \vrf/regTable_reg[6][95]  ( .E(n3585), .D(\vrf/N113 ), .Q(
        \vrf/regTable[6][95] ) );
  LHQD1BWP \vrf/regTable_reg[6][96]  ( .E(n3585), .D(\vrf/N114 ), .Q(
        \vrf/regTable[6][96] ) );
  LHQD1BWP \vrf/regTable_reg[6][97]  ( .E(n3585), .D(\vrf/N115 ), .Q(
        \vrf/regTable[6][97] ) );
  LHQD1BWP \vrf/regTable_reg[6][98]  ( .E(n3585), .D(\vrf/N116 ), .Q(
        \vrf/regTable[6][98] ) );
  LHQD1BWP \vrf/regTable_reg[6][99]  ( .E(n3585), .D(\vrf/N118 ), .Q(
        \vrf/regTable[6][99] ) );
  LHQD1BWP \vrf/regTable_reg[6][100]  ( .E(n3585), .D(\vrf/N119 ), .Q(
        \vrf/regTable[6][100] ) );
  LHQD1BWP \vrf/regTable_reg[6][101]  ( .E(n3585), .D(\vrf/N120 ), .Q(
        \vrf/regTable[6][101] ) );
  LHQD1BWP \vrf/regTable_reg[6][102]  ( .E(n3585), .D(\vrf/N121 ), .Q(
        \vrf/regTable[6][102] ) );
  LHQD1BWP \vrf/regTable_reg[6][103]  ( .E(n3585), .D(\vrf/N122 ), .Q(
        \vrf/regTable[6][103] ) );
  LHQD1BWP \vrf/regTable_reg[6][104]  ( .E(n3585), .D(\vrf/N123 ), .Q(
        \vrf/regTable[6][104] ) );
  LHQD1BWP \vrf/regTable_reg[6][105]  ( .E(n3585), .D(\vrf/N124 ), .Q(
        \vrf/regTable[6][105] ) );
  LHQD1BWP \vrf/regTable_reg[6][106]  ( .E(n3585), .D(\vrf/N125 ), .Q(
        \vrf/regTable[6][106] ) );
  LHQD1BWP \vrf/regTable_reg[6][107]  ( .E(n3585), .D(\vrf/N126 ), .Q(
        \vrf/regTable[6][107] ) );
  LHQD1BWP \vrf/regTable_reg[6][108]  ( .E(n3585), .D(\vrf/N127 ), .Q(
        \vrf/regTable[6][108] ) );
  LHQD1BWP \vrf/regTable_reg[6][109]  ( .E(n3585), .D(\vrf/N128 ), .Q(
        \vrf/regTable[6][109] ) );
  LHQD1BWP \vrf/regTable_reg[6][110]  ( .E(n3585), .D(\vrf/N129 ), .Q(
        \vrf/regTable[6][110] ) );
  LHQD1BWP \vrf/regTable_reg[6][111]  ( .E(n3585), .D(\vrf/N130 ), .Q(
        \vrf/regTable[6][111] ) );
  LHQD1BWP \vrf/regTable_reg[6][112]  ( .E(n3585), .D(\vrf/N131 ), .Q(
        \vrf/regTable[6][112] ) );
  LHQD1BWP \vrf/regTable_reg[6][113]  ( .E(n3585), .D(\vrf/N132 ), .Q(
        \vrf/regTable[6][113] ) );
  LHQD1BWP \vrf/regTable_reg[6][114]  ( .E(n3585), .D(\vrf/N133 ), .Q(
        \vrf/regTable[6][114] ) );
  LHQD1BWP \vrf/regTable_reg[6][115]  ( .E(n3585), .D(\vrf/N134 ), .Q(
        \vrf/regTable[6][115] ) );
  LHQD1BWP \vrf/regTable_reg[6][116]  ( .E(n3585), .D(\vrf/N135 ), .Q(
        \vrf/regTable[6][116] ) );
  LHQD1BWP \vrf/regTable_reg[6][117]  ( .E(n3585), .D(\vrf/N136 ), .Q(
        \vrf/regTable[6][117] ) );
  LHQD1BWP \vrf/regTable_reg[6][118]  ( .E(n3585), .D(\vrf/N137 ), .Q(
        \vrf/regTable[6][118] ) );
  LHQD1BWP \vrf/regTable_reg[6][119]  ( .E(n3585), .D(\vrf/N138 ), .Q(
        \vrf/regTable[6][119] ) );
  LHQD1BWP \vrf/regTable_reg[6][120]  ( .E(n3585), .D(\vrf/N139 ), .Q(
        \vrf/regTable[6][120] ) );
  LHQD1BWP \vrf/regTable_reg[6][121]  ( .E(n3585), .D(\vrf/N140 ), .Q(
        \vrf/regTable[6][121] ) );
  LHQD1BWP \vrf/regTable_reg[6][122]  ( .E(n3585), .D(\vrf/N141 ), .Q(
        \vrf/regTable[6][122] ) );
  LHQD1BWP \vrf/regTable_reg[6][123]  ( .E(n3585), .D(\vrf/N142 ), .Q(
        \vrf/regTable[6][123] ) );
  LHQD1BWP \vrf/regTable_reg[6][124]  ( .E(n3585), .D(\vrf/N143 ), .Q(
        \vrf/regTable[6][124] ) );
  LHQD1BWP \vrf/regTable_reg[6][125]  ( .E(n3585), .D(\vrf/N144 ), .Q(
        \vrf/regTable[6][125] ) );
  LHQD1BWP \vrf/regTable_reg[6][126]  ( .E(n3585), .D(\vrf/N145 ), .Q(
        \vrf/regTable[6][126] ) );
  LHQD1BWP \vrf/regTable_reg[6][127]  ( .E(n3585), .D(\vrf/N146 ), .Q(
        \vrf/regTable[6][127] ) );
  LHQD1BWP \vrf/regTable_reg[6][128]  ( .E(n3585), .D(\vrf/N147 ), .Q(
        \vrf/regTable[6][128] ) );
  LHQD1BWP \vrf/regTable_reg[6][129]  ( .E(n3585), .D(\vrf/N148 ), .Q(
        \vrf/regTable[6][129] ) );
  LHQD1BWP \vrf/regTable_reg[6][130]  ( .E(n3585), .D(\vrf/N149 ), .Q(
        \vrf/regTable[6][130] ) );
  LHQD1BWP \vrf/regTable_reg[6][131]  ( .E(n3585), .D(\vrf/N150 ), .Q(
        \vrf/regTable[6][131] ) );
  LHQD1BWP \vrf/regTable_reg[6][132]  ( .E(n3585), .D(\vrf/N151 ), .Q(
        \vrf/regTable[6][132] ) );
  LHQD1BWP \vrf/regTable_reg[6][133]  ( .E(n3585), .D(\vrf/N152 ), .Q(
        \vrf/regTable[6][133] ) );
  LHQD1BWP \vrf/regTable_reg[6][134]  ( .E(n3585), .D(\vrf/N153 ), .Q(
        \vrf/regTable[6][134] ) );
  LHQD1BWP \vrf/regTable_reg[6][135]  ( .E(n3585), .D(\vrf/N154 ), .Q(
        \vrf/regTable[6][135] ) );
  LHQD1BWP \vrf/regTable_reg[6][136]  ( .E(n3585), .D(\vrf/N155 ), .Q(
        \vrf/regTable[6][136] ) );
  LHQD1BWP \vrf/regTable_reg[6][137]  ( .E(\vrf/N278 ), .D(\vrf/N156 ), .Q(
        \vrf/regTable[6][137] ) );
  LHQD1BWP \vrf/regTable_reg[6][138]  ( .E(n3585), .D(\vrf/N157 ), .Q(
        \vrf/regTable[6][138] ) );
  LHQD1BWP \vrf/regTable_reg[6][139]  ( .E(\vrf/N278 ), .D(\vrf/N158 ), .Q(
        \vrf/regTable[6][139] ) );
  LHQD1BWP \vrf/regTable_reg[6][140]  ( .E(n3585), .D(\vrf/N159 ), .Q(
        \vrf/regTable[6][140] ) );
  LHQD1BWP \vrf/regTable_reg[6][141]  ( .E(\vrf/N278 ), .D(\vrf/N160 ), .Q(
        \vrf/regTable[6][141] ) );
  LHQD1BWP \vrf/regTable_reg[6][142]  ( .E(n3585), .D(\vrf/N161 ), .Q(
        \vrf/regTable[6][142] ) );
  LHQD1BWP \vrf/regTable_reg[6][143]  ( .E(\vrf/N278 ), .D(\vrf/N162 ), .Q(
        \vrf/regTable[6][143] ) );
  LHQD1BWP \vrf/regTable_reg[6][144]  ( .E(n3585), .D(\vrf/N163 ), .Q(
        \vrf/regTable[6][144] ) );
  LHQD1BWP \vrf/regTable_reg[6][145]  ( .E(\vrf/N278 ), .D(\vrf/N164 ), .Q(
        \vrf/regTable[6][145] ) );
  LHQD1BWP \vrf/regTable_reg[6][146]  ( .E(n3585), .D(\vrf/N165 ), .Q(
        \vrf/regTable[6][146] ) );
  LHQD1BWP \vrf/regTable_reg[6][147]  ( .E(\vrf/N278 ), .D(\vrf/N166 ), .Q(
        \vrf/regTable[6][147] ) );
  LHQD1BWP \vrf/regTable_reg[6][148]  ( .E(n3585), .D(\vrf/N167 ), .Q(
        \vrf/regTable[6][148] ) );
  LHQD1BWP \vrf/regTable_reg[6][149]  ( .E(n3585), .D(\vrf/N168 ), .Q(
        \vrf/regTable[6][149] ) );
  LHQD1BWP \vrf/regTable_reg[6][150]  ( .E(n3585), .D(\vrf/N169 ), .Q(
        \vrf/regTable[6][150] ) );
  LHQD1BWP \vrf/regTable_reg[6][151]  ( .E(\vrf/N278 ), .D(\vrf/N170 ), .Q(
        \vrf/regTable[6][151] ) );
  LHQD1BWP \vrf/regTable_reg[6][152]  ( .E(n3585), .D(\vrf/N171 ), .Q(
        \vrf/regTable[6][152] ) );
  LHQD1BWP \vrf/regTable_reg[6][153]  ( .E(n3585), .D(\vrf/N172 ), .Q(
        \vrf/regTable[6][153] ) );
  LHQD1BWP \vrf/regTable_reg[6][154]  ( .E(n3585), .D(\vrf/N173 ), .Q(
        \vrf/regTable[6][154] ) );
  LHQD1BWP \vrf/regTable_reg[6][155]  ( .E(\vrf/N278 ), .D(\vrf/N174 ), .Q(
        \vrf/regTable[6][155] ) );
  LHQD1BWP \vrf/regTable_reg[6][156]  ( .E(n3585), .D(\vrf/N175 ), .Q(
        \vrf/regTable[6][156] ) );
  LHQD1BWP \vrf/regTable_reg[6][157]  ( .E(n3585), .D(\vrf/N176 ), .Q(
        \vrf/regTable[6][157] ) );
  LHQD1BWP \vrf/regTable_reg[6][158]  ( .E(n3585), .D(\vrf/N177 ), .Q(
        \vrf/regTable[6][158] ) );
  LHQD1BWP \vrf/regTable_reg[6][159]  ( .E(n3585), .D(\vrf/N178 ), .Q(
        \vrf/regTable[6][159] ) );
  LHQD1BWP \vrf/regTable_reg[6][160]  ( .E(\vrf/N278 ), .D(\vrf/N179 ), .Q(
        \vrf/regTable[6][160] ) );
  LHQD1BWP \vrf/regTable_reg[6][161]  ( .E(n3585), .D(\vrf/N180 ), .Q(
        \vrf/regTable[6][161] ) );
  LHQD1BWP \vrf/regTable_reg[6][162]  ( .E(n3585), .D(\vrf/N181 ), .Q(
        \vrf/regTable[6][162] ) );
  LHQD1BWP \vrf/regTable_reg[6][163]  ( .E(n3585), .D(\vrf/N182 ), .Q(
        \vrf/regTable[6][163] ) );
  LHQD1BWP \vrf/regTable_reg[6][164]  ( .E(\vrf/N278 ), .D(\vrf/N183 ), .Q(
        \vrf/regTable[6][164] ) );
  LHQD1BWP \vrf/regTable_reg[6][165]  ( .E(n3585), .D(\vrf/N184 ), .Q(
        \vrf/regTable[6][165] ) );
  LHQD1BWP \vrf/regTable_reg[6][166]  ( .E(n3585), .D(\vrf/N185 ), .Q(
        \vrf/regTable[6][166] ) );
  LHQD1BWP \vrf/regTable_reg[6][167]  ( .E(n3585), .D(\vrf/N186 ), .Q(
        \vrf/regTable[6][167] ) );
  LHQD1BWP \vrf/regTable_reg[6][168]  ( .E(\vrf/N278 ), .D(\vrf/N187 ), .Q(
        \vrf/regTable[6][168] ) );
  LHQD1BWP \vrf/regTable_reg[6][169]  ( .E(n3585), .D(\vrf/N188 ), .Q(
        \vrf/regTable[6][169] ) );
  LHQD1BWP \vrf/regTable_reg[6][170]  ( .E(n3585), .D(\vrf/N189 ), .Q(
        \vrf/regTable[6][170] ) );
  LHQD1BWP \vrf/regTable_reg[6][171]  ( .E(n3585), .D(\vrf/N190 ), .Q(
        \vrf/regTable[6][171] ) );
  LHQD1BWP \vrf/regTable_reg[6][172]  ( .E(n3585), .D(\vrf/N191 ), .Q(
        \vrf/regTable[6][172] ) );
  LHQD1BWP \vrf/regTable_reg[6][173]  ( .E(n3585), .D(\vrf/N192 ), .Q(
        \vrf/regTable[6][173] ) );
  LHQD1BWP \vrf/regTable_reg[6][174]  ( .E(\vrf/N278 ), .D(\vrf/N193 ), .Q(
        \vrf/regTable[6][174] ) );
  LHQD1BWP \vrf/regTable_reg[6][175]  ( .E(n3585), .D(\vrf/N194 ), .Q(
        \vrf/regTable[6][175] ) );
  LHQD1BWP \vrf/regTable_reg[6][176]  ( .E(n3585), .D(\vrf/N195 ), .Q(
        \vrf/regTable[6][176] ) );
  LHQD1BWP \vrf/regTable_reg[6][177]  ( .E(n3585), .D(\vrf/N196 ), .Q(
        \vrf/regTable[6][177] ) );
  LHQD1BWP \vrf/regTable_reg[6][178]  ( .E(n3585), .D(\vrf/N197 ), .Q(
        \vrf/regTable[6][178] ) );
  LHQD1BWP \vrf/regTable_reg[6][179]  ( .E(\vrf/N278 ), .D(\vrf/N198 ), .Q(
        \vrf/regTable[6][179] ) );
  LHQD1BWP \vrf/regTable_reg[6][180]  ( .E(n3585), .D(\vrf/N199 ), .Q(
        \vrf/regTable[6][180] ) );
  LHQD1BWP \vrf/regTable_reg[6][181]  ( .E(n3585), .D(\vrf/N200 ), .Q(
        \vrf/regTable[6][181] ) );
  LHQD1BWP \vrf/regTable_reg[6][182]  ( .E(n3585), .D(\vrf/N201 ), .Q(
        \vrf/regTable[6][182] ) );
  LHQD1BWP \vrf/regTable_reg[6][183]  ( .E(n3585), .D(\vrf/N202 ), .Q(
        \vrf/regTable[6][183] ) );
  LHQD1BWP \vrf/regTable_reg[6][184]  ( .E(n3585), .D(\vrf/N203 ), .Q(
        \vrf/regTable[6][184] ) );
  LHQD1BWP \vrf/regTable_reg[6][185]  ( .E(n3585), .D(\vrf/N204 ), .Q(
        \vrf/regTable[6][185] ) );
  LHQD1BWP \vrf/regTable_reg[6][186]  ( .E(n3585), .D(\vrf/N205 ), .Q(
        \vrf/regTable[6][186] ) );
  LHQD1BWP \vrf/regTable_reg[6][187]  ( .E(n3585), .D(\vrf/N206 ), .Q(
        \vrf/regTable[6][187] ) );
  LHQD1BWP \vrf/regTable_reg[6][188]  ( .E(n3585), .D(\vrf/N207 ), .Q(
        \vrf/regTable[6][188] ) );
  LHQD1BWP \vrf/regTable_reg[6][189]  ( .E(\vrf/N278 ), .D(\vrf/N208 ), .Q(
        \vrf/regTable[6][189] ) );
  LHQD1BWP \vrf/regTable_reg[6][190]  ( .E(n3585), .D(\vrf/N209 ), .Q(
        \vrf/regTable[6][190] ) );
  LHQD1BWP \vrf/regTable_reg[6][191]  ( .E(n3585), .D(\vrf/N210 ), .Q(
        \vrf/regTable[6][191] ) );
  LHQD1BWP \vrf/regTable_reg[6][192]  ( .E(n3585), .D(\vrf/N211 ), .Q(
        \vrf/regTable[6][192] ) );
  LHQD1BWP \vrf/regTable_reg[6][193]  ( .E(n3585), .D(\vrf/N212 ), .Q(
        \vrf/regTable[6][193] ) );
  LHQD1BWP \vrf/regTable_reg[6][194]  ( .E(\vrf/N278 ), .D(\vrf/N213 ), .Q(
        \vrf/regTable[6][194] ) );
  LHQD1BWP \vrf/regTable_reg[6][195]  ( .E(\vrf/N278 ), .D(\vrf/N214 ), .Q(
        \vrf/regTable[6][195] ) );
  LHQD1BWP \vrf/regTable_reg[6][196]  ( .E(n3585), .D(\vrf/N215 ), .Q(
        \vrf/regTable[6][196] ) );
  LHQD1BWP \vrf/regTable_reg[6][197]  ( .E(n3585), .D(\vrf/N216 ), .Q(
        \vrf/regTable[6][197] ) );
  LHQD1BWP \vrf/regTable_reg[6][198]  ( .E(n3585), .D(\vrf/N218 ), .Q(
        \vrf/regTable[6][198] ) );
  LHQD1BWP \vrf/regTable_reg[6][199]  ( .E(n3585), .D(\vrf/N219 ), .Q(
        \vrf/regTable[6][199] ) );
  LHQD1BWP \vrf/regTable_reg[6][200]  ( .E(n3585), .D(\vrf/N220 ), .Q(
        \vrf/regTable[6][200] ) );
  LHQD1BWP \vrf/regTable_reg[6][201]  ( .E(\vrf/N278 ), .D(\vrf/N221 ), .Q(
        \vrf/regTable[6][201] ) );
  LHQD1BWP \vrf/regTable_reg[6][202]  ( .E(n3585), .D(\vrf/N222 ), .Q(
        \vrf/regTable[6][202] ) );
  LHQD1BWP \vrf/regTable_reg[6][203]  ( .E(n3585), .D(\vrf/N223 ), .Q(
        \vrf/regTable[6][203] ) );
  LHQD1BWP \vrf/regTable_reg[6][204]  ( .E(\vrf/N278 ), .D(\vrf/N224 ), .Q(
        \vrf/regTable[6][204] ) );
  LHQD1BWP \vrf/regTable_reg[6][205]  ( .E(n3585), .D(\vrf/N225 ), .Q(
        \vrf/regTable[6][205] ) );
  LHQD1BWP \vrf/regTable_reg[6][206]  ( .E(\vrf/N278 ), .D(\vrf/N226 ), .Q(
        \vrf/regTable[6][206] ) );
  LHQD1BWP \vrf/regTable_reg[6][207]  ( .E(n3585), .D(\vrf/N227 ), .Q(
        \vrf/regTable[6][207] ) );
  LHQD1BWP \vrf/regTable_reg[6][208]  ( .E(n3585), .D(\vrf/N228 ), .Q(
        \vrf/regTable[6][208] ) );
  LHQD1BWP \vrf/regTable_reg[6][209]  ( .E(n3585), .D(\vrf/N229 ), .Q(
        \vrf/regTable[6][209] ) );
  LHQD1BWP \vrf/regTable_reg[6][210]  ( .E(n3585), .D(\vrf/N230 ), .Q(
        \vrf/regTable[6][210] ) );
  LHQD1BWP \vrf/regTable_reg[6][211]  ( .E(n3585), .D(\vrf/N231 ), .Q(
        \vrf/regTable[6][211] ) );
  LHQD1BWP \vrf/regTable_reg[6][212]  ( .E(n3585), .D(\vrf/N232 ), .Q(
        \vrf/regTable[6][212] ) );
  LHQD1BWP \vrf/regTable_reg[6][213]  ( .E(n3585), .D(\vrf/N233 ), .Q(
        \vrf/regTable[6][213] ) );
  LHQD1BWP \vrf/regTable_reg[6][214]  ( .E(n3585), .D(\vrf/N234 ), .Q(
        \vrf/regTable[6][214] ) );
  LHQD1BWP \vrf/regTable_reg[6][215]  ( .E(n3585), .D(\vrf/N235 ), .Q(
        \vrf/regTable[6][215] ) );
  LHQD1BWP \vrf/regTable_reg[6][216]  ( .E(n3585), .D(\vrf/N236 ), .Q(
        \vrf/regTable[6][216] ) );
  LHQD1BWP \vrf/regTable_reg[6][217]  ( .E(n3585), .D(\vrf/N237 ), .Q(
        \vrf/regTable[6][217] ) );
  LHQD1BWP \vrf/regTable_reg[6][218]  ( .E(n3585), .D(\vrf/N238 ), .Q(
        \vrf/regTable[6][218] ) );
  LHQD1BWP \vrf/regTable_reg[6][219]  ( .E(n3585), .D(\vrf/N239 ), .Q(
        \vrf/regTable[6][219] ) );
  LHQD1BWP \vrf/regTable_reg[6][220]  ( .E(n3585), .D(\vrf/N240 ), .Q(
        \vrf/regTable[6][220] ) );
  LHQD1BWP \vrf/regTable_reg[6][221]  ( .E(n3585), .D(\vrf/N241 ), .Q(
        \vrf/regTable[6][221] ) );
  LHQD1BWP \vrf/regTable_reg[6][222]  ( .E(n3585), .D(\vrf/N242 ), .Q(
        \vrf/regTable[6][222] ) );
  LHQD1BWP \vrf/regTable_reg[6][223]  ( .E(\vrf/N278 ), .D(\vrf/N243 ), .Q(
        \vrf/regTable[6][223] ) );
  LHQD1BWP \vrf/regTable_reg[6][224]  ( .E(n3585), .D(\vrf/N244 ), .Q(
        \vrf/regTable[6][224] ) );
  LHQD1BWP \vrf/regTable_reg[6][225]  ( .E(n3585), .D(\vrf/N245 ), .Q(
        \vrf/regTable[6][225] ) );
  LHQD1BWP \vrf/regTable_reg[6][226]  ( .E(n3585), .D(\vrf/N246 ), .Q(
        \vrf/regTable[6][226] ) );
  LHQD1BWP \vrf/regTable_reg[6][227]  ( .E(\vrf/N278 ), .D(\vrf/N247 ), .Q(
        \vrf/regTable[6][227] ) );
  LHQD1BWP \vrf/regTable_reg[6][228]  ( .E(n3585), .D(\vrf/N248 ), .Q(
        \vrf/regTable[6][228] ) );
  LHQD1BWP \vrf/regTable_reg[6][229]  ( .E(n3585), .D(\vrf/N249 ), .Q(
        \vrf/regTable[6][229] ) );
  LHQD1BWP \vrf/regTable_reg[6][230]  ( .E(n3585), .D(\vrf/N250 ), .Q(
        \vrf/regTable[6][230] ) );
  LHQD1BWP \vrf/regTable_reg[6][231]  ( .E(\vrf/N278 ), .D(\vrf/N251 ), .Q(
        \vrf/regTable[6][231] ) );
  LHQD1BWP \vrf/regTable_reg[6][232]  ( .E(n3585), .D(\vrf/N252 ), .Q(
        \vrf/regTable[6][232] ) );
  LHQD1BWP \vrf/regTable_reg[6][233]  ( .E(n3585), .D(\vrf/N253 ), .Q(
        \vrf/regTable[6][233] ) );
  LHQD1BWP \vrf/regTable_reg[6][234]  ( .E(n3585), .D(\vrf/N254 ), .Q(
        \vrf/regTable[6][234] ) );
  LHQD1BWP \vrf/regTable_reg[6][235]  ( .E(n3585), .D(\vrf/N255 ), .Q(
        \vrf/regTable[6][235] ) );
  LHQD1BWP \vrf/regTable_reg[6][236]  ( .E(n3585), .D(\vrf/N256 ), .Q(
        \vrf/regTable[6][236] ) );
  LHQD1BWP \vrf/regTable_reg[6][237]  ( .E(n3585), .D(\vrf/N257 ), .Q(
        \vrf/regTable[6][237] ) );
  LHQD1BWP \vrf/regTable_reg[6][238]  ( .E(n3585), .D(\vrf/N258 ), .Q(
        \vrf/regTable[6][238] ) );
  LHQD1BWP \vrf/regTable_reg[6][239]  ( .E(n3585), .D(\vrf/N259 ), .Q(
        \vrf/regTable[6][239] ) );
  LHQD1BWP \vrf/regTable_reg[6][240]  ( .E(n3585), .D(\vrf/N260 ), .Q(
        \vrf/regTable[6][240] ) );
  LHQD1BWP \vrf/regTable_reg[6][241]  ( .E(n3585), .D(\vrf/N261 ), .Q(
        \vrf/regTable[6][241] ) );
  LHQD1BWP \vrf/regTable_reg[6][242]  ( .E(n3585), .D(\vrf/N262 ), .Q(
        \vrf/regTable[6][242] ) );
  LHQD1BWP \vrf/regTable_reg[6][243]  ( .E(n3585), .D(\vrf/N263 ), .Q(
        \vrf/regTable[6][243] ) );
  LHQD1BWP \vrf/regTable_reg[6][244]  ( .E(n3585), .D(\vrf/N264 ), .Q(
        \vrf/regTable[6][244] ) );
  LHQD1BWP \vrf/regTable_reg[6][245]  ( .E(n3585), .D(\vrf/N265 ), .Q(
        \vrf/regTable[6][245] ) );
  LHQD1BWP \vrf/regTable_reg[6][246]  ( .E(n3585), .D(\vrf/N266 ), .Q(
        \vrf/regTable[6][246] ) );
  LHQD1BWP \vrf/regTable_reg[6][247]  ( .E(n3585), .D(\vrf/N267 ), .Q(
        \vrf/regTable[6][247] ) );
  LHQD1BWP \vrf/regTable_reg[6][248]  ( .E(n3585), .D(\vrf/N268 ), .Q(
        \vrf/regTable[6][248] ) );
  LHQD1BWP \vrf/regTable_reg[6][249]  ( .E(n3585), .D(\vrf/N269 ), .Q(
        \vrf/regTable[6][249] ) );
  LHQD1BWP \vrf/regTable_reg[6][250]  ( .E(n3585), .D(\vrf/N270 ), .Q(
        \vrf/regTable[6][250] ) );
  LHQD1BWP \vrf/regTable_reg[6][251]  ( .E(\vrf/N278 ), .D(\vrf/N271 ), .Q(
        \vrf/regTable[6][251] ) );
  LHQD1BWP \vrf/regTable_reg[6][252]  ( .E(n3585), .D(\vrf/N272 ), .Q(
        \vrf/regTable[6][252] ) );
  LHQD1BWP \vrf/regTable_reg[6][253]  ( .E(n3585), .D(\vrf/N273 ), .Q(
        \vrf/regTable[6][253] ) );
  LHQD1BWP \vrf/regTable_reg[6][254]  ( .E(n3585), .D(\vrf/N274 ), .Q(
        \vrf/regTable[6][254] ) );
  LHQD1BWP \vrf/regTable_reg[6][255]  ( .E(n3585), .D(\vrf/N275 ), .Q(
        \vrf/regTable[6][255] ) );
  LHQD1BWP \vrf/regTable_reg[5][0]  ( .E(n3584), .D(\vrf/N18 ), .Q(
        \vrf/regTable[5][0] ) );
  LHQD1BWP \vrf/regTable_reg[5][1]  ( .E(n3584), .D(\vrf/N19 ), .Q(
        \vrf/regTable[5][1] ) );
  LHQD1BWP \vrf/regTable_reg[5][2]  ( .E(n3584), .D(\vrf/N20 ), .Q(
        \vrf/regTable[5][2] ) );
  LHQD1BWP \vrf/regTable_reg[5][3]  ( .E(n3584), .D(\vrf/N21 ), .Q(
        \vrf/regTable[5][3] ) );
  LHQD1BWP \vrf/regTable_reg[5][4]  ( .E(n3584), .D(\vrf/N22 ), .Q(
        \vrf/regTable[5][4] ) );
  LHQD1BWP \vrf/regTable_reg[5][5]  ( .E(n3584), .D(\vrf/N23 ), .Q(
        \vrf/regTable[5][5] ) );
  LHQD1BWP \vrf/regTable_reg[5][6]  ( .E(n3584), .D(\vrf/N24 ), .Q(
        \vrf/regTable[5][6] ) );
  LHQD1BWP \vrf/regTable_reg[5][7]  ( .E(n3584), .D(\vrf/N25 ), .Q(
        \vrf/regTable[5][7] ) );
  LHQD1BWP \vrf/regTable_reg[5][8]  ( .E(n3584), .D(\vrf/N26 ), .Q(
        \vrf/regTable[5][8] ) );
  LHQD1BWP \vrf/regTable_reg[5][9]  ( .E(n3584), .D(\vrf/N27 ), .Q(
        \vrf/regTable[5][9] ) );
  LHQD1BWP \vrf/regTable_reg[5][10]  ( .E(n3584), .D(\vrf/N28 ), .Q(
        \vrf/regTable[5][10] ) );
  LHQD1BWP \vrf/regTable_reg[5][11]  ( .E(n3584), .D(\vrf/N29 ), .Q(
        \vrf/regTable[5][11] ) );
  LHQD1BWP \vrf/regTable_reg[5][12]  ( .E(n3584), .D(\vrf/N30 ), .Q(
        \vrf/regTable[5][12] ) );
  LHQD1BWP \vrf/regTable_reg[5][13]  ( .E(n3584), .D(\vrf/N31 ), .Q(
        \vrf/regTable[5][13] ) );
  LHQD1BWP \vrf/regTable_reg[5][14]  ( .E(n3584), .D(\vrf/N32 ), .Q(
        \vrf/regTable[5][14] ) );
  LHQD1BWP \vrf/regTable_reg[5][15]  ( .E(n3584), .D(\vrf/N33 ), .Q(
        \vrf/regTable[5][15] ) );
  LHQD1BWP \vrf/regTable_reg[5][16]  ( .E(n3584), .D(\vrf/N34 ), .Q(
        \vrf/regTable[5][16] ) );
  LHQD1BWP \vrf/regTable_reg[5][17]  ( .E(n3584), .D(\vrf/N35 ), .Q(
        \vrf/regTable[5][17] ) );
  LHQD1BWP \vrf/regTable_reg[5][18]  ( .E(n3584), .D(\vrf/N36 ), .Q(
        \vrf/regTable[5][18] ) );
  LHQD1BWP \vrf/regTable_reg[5][19]  ( .E(n3584), .D(\vrf/N37 ), .Q(
        \vrf/regTable[5][19] ) );
  LHQD1BWP \vrf/regTable_reg[5][20]  ( .E(n3584), .D(\vrf/N38 ), .Q(
        \vrf/regTable[5][20] ) );
  LHQD1BWP \vrf/regTable_reg[5][21]  ( .E(n3584), .D(\vrf/N39 ), .Q(
        \vrf/regTable[5][21] ) );
  LHQD1BWP \vrf/regTable_reg[5][22]  ( .E(n3584), .D(\vrf/N40 ), .Q(
        \vrf/regTable[5][22] ) );
  LHQD1BWP \vrf/regTable_reg[5][23]  ( .E(n3584), .D(\vrf/N41 ), .Q(
        \vrf/regTable[5][23] ) );
  LHQD1BWP \vrf/regTable_reg[5][24]  ( .E(n3584), .D(\vrf/N42 ), .Q(
        \vrf/regTable[5][24] ) );
  LHQD1BWP \vrf/regTable_reg[5][25]  ( .E(n3584), .D(\vrf/N43 ), .Q(
        \vrf/regTable[5][25] ) );
  LHQD1BWP \vrf/regTable_reg[5][26]  ( .E(n3584), .D(\vrf/N44 ), .Q(
        \vrf/regTable[5][26] ) );
  LHQD1BWP \vrf/regTable_reg[5][27]  ( .E(n3584), .D(\vrf/N45 ), .Q(
        \vrf/regTable[5][27] ) );
  LHQD1BWP \vrf/regTable_reg[5][28]  ( .E(n3584), .D(\vrf/N46 ), .Q(
        \vrf/regTable[5][28] ) );
  LHQD1BWP \vrf/regTable_reg[5][29]  ( .E(n3584), .D(\vrf/N47 ), .Q(
        \vrf/regTable[5][29] ) );
  LHQD1BWP \vrf/regTable_reg[5][30]  ( .E(n3584), .D(\vrf/N48 ), .Q(
        \vrf/regTable[5][30] ) );
  LHQD1BWP \vrf/regTable_reg[5][31]  ( .E(n3584), .D(\vrf/N49 ), .Q(
        \vrf/regTable[5][31] ) );
  LHQD1BWP \vrf/regTable_reg[5][32]  ( .E(n3584), .D(\vrf/N50 ), .Q(
        \vrf/regTable[5][32] ) );
  LHQD1BWP \vrf/regTable_reg[5][33]  ( .E(n3584), .D(\vrf/N51 ), .Q(
        \vrf/regTable[5][33] ) );
  LHQD1BWP \vrf/regTable_reg[5][34]  ( .E(n3584), .D(\vrf/N52 ), .Q(
        \vrf/regTable[5][34] ) );
  LHQD1BWP \vrf/regTable_reg[5][35]  ( .E(n3584), .D(\vrf/N53 ), .Q(
        \vrf/regTable[5][35] ) );
  LHQD1BWP \vrf/regTable_reg[5][36]  ( .E(n3584), .D(\vrf/N54 ), .Q(
        \vrf/regTable[5][36] ) );
  LHQD1BWP \vrf/regTable_reg[5][37]  ( .E(n3584), .D(\vrf/N55 ), .Q(
        \vrf/regTable[5][37] ) );
  LHQD1BWP \vrf/regTable_reg[5][38]  ( .E(n3584), .D(\vrf/N56 ), .Q(
        \vrf/regTable[5][38] ) );
  LHQD1BWP \vrf/regTable_reg[5][39]  ( .E(n3584), .D(\vrf/N57 ), .Q(
        \vrf/regTable[5][39] ) );
  LHQD1BWP \vrf/regTable_reg[5][40]  ( .E(n3584), .D(\vrf/N58 ), .Q(
        \vrf/regTable[5][40] ) );
  LHQD1BWP \vrf/regTable_reg[5][41]  ( .E(n3584), .D(\vrf/N59 ), .Q(
        \vrf/regTable[5][41] ) );
  LHQD1BWP \vrf/regTable_reg[5][42]  ( .E(n3584), .D(\vrf/N60 ), .Q(
        \vrf/regTable[5][42] ) );
  LHQD1BWP \vrf/regTable_reg[5][43]  ( .E(n3584), .D(\vrf/N61 ), .Q(
        \vrf/regTable[5][43] ) );
  LHQD1BWP \vrf/regTable_reg[5][44]  ( .E(n3584), .D(\vrf/N62 ), .Q(
        \vrf/regTable[5][44] ) );
  LHQD1BWP \vrf/regTable_reg[5][45]  ( .E(n3584), .D(\vrf/N63 ), .Q(
        \vrf/regTable[5][45] ) );
  LHQD1BWP \vrf/regTable_reg[5][46]  ( .E(n3584), .D(\vrf/N64 ), .Q(
        \vrf/regTable[5][46] ) );
  LHQD1BWP \vrf/regTable_reg[5][47]  ( .E(n3584), .D(\vrf/N65 ), .Q(
        \vrf/regTable[5][47] ) );
  LHQD1BWP \vrf/regTable_reg[5][48]  ( .E(n3584), .D(\vrf/N66 ), .Q(
        \vrf/regTable[5][48] ) );
  LHQD1BWP \vrf/regTable_reg[5][49]  ( .E(n3584), .D(\vrf/N67 ), .Q(
        \vrf/regTable[5][49] ) );
  LHQD1BWP \vrf/regTable_reg[5][50]  ( .E(n3584), .D(\vrf/N68 ), .Q(
        \vrf/regTable[5][50] ) );
  LHQD1BWP \vrf/regTable_reg[5][51]  ( .E(n3584), .D(\vrf/N69 ), .Q(
        \vrf/regTable[5][51] ) );
  LHQD1BWP \vrf/regTable_reg[5][52]  ( .E(n3584), .D(\vrf/N70 ), .Q(
        \vrf/regTable[5][52] ) );
  LHQD1BWP \vrf/regTable_reg[5][53]  ( .E(n3584), .D(\vrf/N71 ), .Q(
        \vrf/regTable[5][53] ) );
  LHQD1BWP \vrf/regTable_reg[5][54]  ( .E(n3584), .D(\vrf/N72 ), .Q(
        \vrf/regTable[5][54] ) );
  LHQD1BWP \vrf/regTable_reg[5][55]  ( .E(n3584), .D(\vrf/N73 ), .Q(
        \vrf/regTable[5][55] ) );
  LHQD1BWP \vrf/regTable_reg[5][56]  ( .E(n3584), .D(\vrf/N74 ), .Q(
        \vrf/regTable[5][56] ) );
  LHQD1BWP \vrf/regTable_reg[5][57]  ( .E(n3584), .D(\vrf/N75 ), .Q(
        \vrf/regTable[5][57] ) );
  LHQD1BWP \vrf/regTable_reg[5][58]  ( .E(n3584), .D(\vrf/N76 ), .Q(
        \vrf/regTable[5][58] ) );
  LHQD1BWP \vrf/regTable_reg[5][59]  ( .E(n3584), .D(\vrf/N77 ), .Q(
        \vrf/regTable[5][59] ) );
  LHQD1BWP \vrf/regTable_reg[5][60]  ( .E(n3584), .D(\vrf/N78 ), .Q(
        \vrf/regTable[5][60] ) );
  LHQD1BWP \vrf/regTable_reg[5][61]  ( .E(n3584), .D(\vrf/N79 ), .Q(
        \vrf/regTable[5][61] ) );
  LHQD1BWP \vrf/regTable_reg[5][62]  ( .E(n3584), .D(\vrf/N80 ), .Q(
        \vrf/regTable[5][62] ) );
  LHQD1BWP \vrf/regTable_reg[5][63]  ( .E(n3584), .D(\vrf/N81 ), .Q(
        \vrf/regTable[5][63] ) );
  LHQD1BWP \vrf/regTable_reg[5][64]  ( .E(n3584), .D(\vrf/N82 ), .Q(
        \vrf/regTable[5][64] ) );
  LHQD1BWP \vrf/regTable_reg[5][65]  ( .E(n3584), .D(\vrf/N83 ), .Q(
        \vrf/regTable[5][65] ) );
  LHQD1BWP \vrf/regTable_reg[5][66]  ( .E(n3584), .D(\vrf/N84 ), .Q(
        \vrf/regTable[5][66] ) );
  LHQD1BWP \vrf/regTable_reg[5][67]  ( .E(n3584), .D(\vrf/N85 ), .Q(
        \vrf/regTable[5][67] ) );
  LHQD1BWP \vrf/regTable_reg[5][68]  ( .E(n3584), .D(\vrf/N86 ), .Q(
        \vrf/regTable[5][68] ) );
  LHQD1BWP \vrf/regTable_reg[5][69]  ( .E(n3584), .D(\vrf/N87 ), .Q(
        \vrf/regTable[5][69] ) );
  LHQD1BWP \vrf/regTable_reg[5][70]  ( .E(n3584), .D(\vrf/N88 ), .Q(
        \vrf/regTable[5][70] ) );
  LHQD1BWP \vrf/regTable_reg[5][71]  ( .E(n3584), .D(\vrf/N89 ), .Q(
        \vrf/regTable[5][71] ) );
  LHQD1BWP \vrf/regTable_reg[5][72]  ( .E(n3584), .D(\vrf/N90 ), .Q(
        \vrf/regTable[5][72] ) );
  LHQD1BWP \vrf/regTable_reg[5][73]  ( .E(n3584), .D(\vrf/N91 ), .Q(
        \vrf/regTable[5][73] ) );
  LHQD1BWP \vrf/regTable_reg[5][74]  ( .E(n3584), .D(\vrf/N92 ), .Q(
        \vrf/regTable[5][74] ) );
  LHQD1BWP \vrf/regTable_reg[5][75]  ( .E(n3584), .D(\vrf/N93 ), .Q(
        \vrf/regTable[5][75] ) );
  LHQD1BWP \vrf/regTable_reg[5][76]  ( .E(n3584), .D(\vrf/N94 ), .Q(
        \vrf/regTable[5][76] ) );
  LHQD1BWP \vrf/regTable_reg[5][77]  ( .E(n3584), .D(\vrf/N95 ), .Q(
        \vrf/regTable[5][77] ) );
  LHQD1BWP \vrf/regTable_reg[5][78]  ( .E(n3584), .D(\vrf/N96 ), .Q(
        \vrf/regTable[5][78] ) );
  LHQD1BWP \vrf/regTable_reg[5][79]  ( .E(n3584), .D(\vrf/N97 ), .Q(
        \vrf/regTable[5][79] ) );
  LHQD1BWP \vrf/regTable_reg[5][80]  ( .E(n3584), .D(\vrf/N98 ), .Q(
        \vrf/regTable[5][80] ) );
  LHQD1BWP \vrf/regTable_reg[5][81]  ( .E(n3584), .D(\vrf/N99 ), .Q(
        \vrf/regTable[5][81] ) );
  LHQD1BWP \vrf/regTable_reg[5][82]  ( .E(n3584), .D(\vrf/N100 ), .Q(
        \vrf/regTable[5][82] ) );
  LHQD1BWP \vrf/regTable_reg[5][83]  ( .E(n3584), .D(\vrf/N101 ), .Q(
        \vrf/regTable[5][83] ) );
  LHQD1BWP \vrf/regTable_reg[5][84]  ( .E(n3584), .D(\vrf/N102 ), .Q(
        \vrf/regTable[5][84] ) );
  LHQD1BWP \vrf/regTable_reg[5][85]  ( .E(n3584), .D(\vrf/N103 ), .Q(
        \vrf/regTable[5][85] ) );
  LHQD1BWP \vrf/regTable_reg[5][86]  ( .E(n3584), .D(\vrf/N104 ), .Q(
        \vrf/regTable[5][86] ) );
  LHQD1BWP \vrf/regTable_reg[5][87]  ( .E(n3584), .D(\vrf/N105 ), .Q(
        \vrf/regTable[5][87] ) );
  LHQD1BWP \vrf/regTable_reg[5][88]  ( .E(n3584), .D(\vrf/N106 ), .Q(
        \vrf/regTable[5][88] ) );
  LHQD1BWP \vrf/regTable_reg[5][89]  ( .E(n3584), .D(\vrf/N107 ), .Q(
        \vrf/regTable[5][89] ) );
  LHQD1BWP \vrf/regTable_reg[5][90]  ( .E(n3584), .D(\vrf/N108 ), .Q(
        \vrf/regTable[5][90] ) );
  LHQD1BWP \vrf/regTable_reg[5][91]  ( .E(n3584), .D(\vrf/N109 ), .Q(
        \vrf/regTable[5][91] ) );
  LHQD1BWP \vrf/regTable_reg[5][92]  ( .E(n3584), .D(\vrf/N110 ), .Q(
        \vrf/regTable[5][92] ) );
  LHQD1BWP \vrf/regTable_reg[5][93]  ( .E(n3584), .D(\vrf/N111 ), .Q(
        \vrf/regTable[5][93] ) );
  LHQD1BWP \vrf/regTable_reg[5][94]  ( .E(n3584), .D(\vrf/N112 ), .Q(
        \vrf/regTable[5][94] ) );
  LHQD1BWP \vrf/regTable_reg[5][95]  ( .E(n3584), .D(\vrf/N113 ), .Q(
        \vrf/regTable[5][95] ) );
  LHQD1BWP \vrf/regTable_reg[5][96]  ( .E(n3584), .D(\vrf/N114 ), .Q(
        \vrf/regTable[5][96] ) );
  LHQD1BWP \vrf/regTable_reg[5][97]  ( .E(n3584), .D(\vrf/N115 ), .Q(
        \vrf/regTable[5][97] ) );
  LHQD1BWP \vrf/regTable_reg[5][98]  ( .E(n3584), .D(\vrf/N116 ), .Q(
        \vrf/regTable[5][98] ) );
  LHQD1BWP \vrf/regTable_reg[5][99]  ( .E(n3584), .D(\vrf/N118 ), .Q(
        \vrf/regTable[5][99] ) );
  LHQD1BWP \vrf/regTable_reg[5][100]  ( .E(n3584), .D(\vrf/N119 ), .Q(
        \vrf/regTable[5][100] ) );
  LHQD1BWP \vrf/regTable_reg[5][101]  ( .E(n3584), .D(\vrf/N120 ), .Q(
        \vrf/regTable[5][101] ) );
  LHQD1BWP \vrf/regTable_reg[5][102]  ( .E(n3584), .D(\vrf/N121 ), .Q(
        \vrf/regTable[5][102] ) );
  LHQD1BWP \vrf/regTable_reg[5][103]  ( .E(n3584), .D(\vrf/N122 ), .Q(
        \vrf/regTable[5][103] ) );
  LHQD1BWP \vrf/regTable_reg[5][104]  ( .E(n3584), .D(\vrf/N123 ), .Q(
        \vrf/regTable[5][104] ) );
  LHQD1BWP \vrf/regTable_reg[5][105]  ( .E(n3584), .D(\vrf/N124 ), .Q(
        \vrf/regTable[5][105] ) );
  LHQD1BWP \vrf/regTable_reg[5][106]  ( .E(n3584), .D(\vrf/N125 ), .Q(
        \vrf/regTable[5][106] ) );
  LHQD1BWP \vrf/regTable_reg[5][107]  ( .E(n3584), .D(\vrf/N126 ), .Q(
        \vrf/regTable[5][107] ) );
  LHQD1BWP \vrf/regTable_reg[5][108]  ( .E(n3584), .D(\vrf/N127 ), .Q(
        \vrf/regTable[5][108] ) );
  LHQD1BWP \vrf/regTable_reg[5][109]  ( .E(n3584), .D(\vrf/N128 ), .Q(
        \vrf/regTable[5][109] ) );
  LHQD1BWP \vrf/regTable_reg[5][110]  ( .E(n3584), .D(\vrf/N129 ), .Q(
        \vrf/regTable[5][110] ) );
  LHQD1BWP \vrf/regTable_reg[5][111]  ( .E(n3584), .D(\vrf/N130 ), .Q(
        \vrf/regTable[5][111] ) );
  LHQD1BWP \vrf/regTable_reg[5][112]  ( .E(n3584), .D(\vrf/N131 ), .Q(
        \vrf/regTable[5][112] ) );
  LHQD1BWP \vrf/regTable_reg[5][113]  ( .E(n3584), .D(\vrf/N132 ), .Q(
        \vrf/regTable[5][113] ) );
  LHQD1BWP \vrf/regTable_reg[5][114]  ( .E(n3584), .D(\vrf/N133 ), .Q(
        \vrf/regTable[5][114] ) );
  LHQD1BWP \vrf/regTable_reg[5][115]  ( .E(n3584), .D(\vrf/N134 ), .Q(
        \vrf/regTable[5][115] ) );
  LHQD1BWP \vrf/regTable_reg[5][116]  ( .E(n3584), .D(\vrf/N135 ), .Q(
        \vrf/regTable[5][116] ) );
  LHQD1BWP \vrf/regTable_reg[5][117]  ( .E(n3584), .D(\vrf/N136 ), .Q(
        \vrf/regTable[5][117] ) );
  LHQD1BWP \vrf/regTable_reg[5][118]  ( .E(n3584), .D(\vrf/N137 ), .Q(
        \vrf/regTable[5][118] ) );
  LHQD1BWP \vrf/regTable_reg[5][119]  ( .E(n3584), .D(\vrf/N138 ), .Q(
        \vrf/regTable[5][119] ) );
  LHQD1BWP \vrf/regTable_reg[5][120]  ( .E(n3584), .D(\vrf/N139 ), .Q(
        \vrf/regTable[5][120] ) );
  LHQD1BWP \vrf/regTable_reg[5][121]  ( .E(n3584), .D(\vrf/N140 ), .Q(
        \vrf/regTable[5][121] ) );
  LHQD1BWP \vrf/regTable_reg[5][122]  ( .E(n3584), .D(\vrf/N141 ), .Q(
        \vrf/regTable[5][122] ) );
  LHQD1BWP \vrf/regTable_reg[5][123]  ( .E(n3584), .D(\vrf/N142 ), .Q(
        \vrf/regTable[5][123] ) );
  LHQD1BWP \vrf/regTable_reg[5][124]  ( .E(n3584), .D(\vrf/N143 ), .Q(
        \vrf/regTable[5][124] ) );
  LHQD1BWP \vrf/regTable_reg[5][125]  ( .E(n3584), .D(\vrf/N144 ), .Q(
        \vrf/regTable[5][125] ) );
  LHQD1BWP \vrf/regTable_reg[5][126]  ( .E(n3584), .D(\vrf/N145 ), .Q(
        \vrf/regTable[5][126] ) );
  LHQD1BWP \vrf/regTable_reg[5][127]  ( .E(n3584), .D(\vrf/N146 ), .Q(
        \vrf/regTable[5][127] ) );
  LHQD1BWP \vrf/regTable_reg[5][128]  ( .E(n3584), .D(\vrf/N147 ), .Q(
        \vrf/regTable[5][128] ) );
  LHQD1BWP \vrf/regTable_reg[5][129]  ( .E(n3584), .D(\vrf/N148 ), .Q(
        \vrf/regTable[5][129] ) );
  LHQD1BWP \vrf/regTable_reg[5][130]  ( .E(n3584), .D(\vrf/N149 ), .Q(
        \vrf/regTable[5][130] ) );
  LHQD1BWP \vrf/regTable_reg[5][131]  ( .E(n3584), .D(\vrf/N150 ), .Q(
        \vrf/regTable[5][131] ) );
  LHQD1BWP \vrf/regTable_reg[5][132]  ( .E(n3584), .D(\vrf/N151 ), .Q(
        \vrf/regTable[5][132] ) );
  LHQD1BWP \vrf/regTable_reg[5][133]  ( .E(n3584), .D(\vrf/N152 ), .Q(
        \vrf/regTable[5][133] ) );
  LHQD1BWP \vrf/regTable_reg[5][134]  ( .E(n3584), .D(\vrf/N153 ), .Q(
        \vrf/regTable[5][134] ) );
  LHQD1BWP \vrf/regTable_reg[5][135]  ( .E(n3584), .D(\vrf/N154 ), .Q(
        \vrf/regTable[5][135] ) );
  LHQD1BWP \vrf/regTable_reg[5][136]  ( .E(n3584), .D(\vrf/N155 ), .Q(
        \vrf/regTable[5][136] ) );
  LHQD1BWP \vrf/regTable_reg[5][137]  ( .E(\vrf/N281 ), .D(\vrf/N156 ), .Q(
        \vrf/regTable[5][137] ) );
  LHQD1BWP \vrf/regTable_reg[5][138]  ( .E(n3584), .D(\vrf/N157 ), .Q(
        \vrf/regTable[5][138] ) );
  LHQD1BWP \vrf/regTable_reg[5][139]  ( .E(\vrf/N281 ), .D(\vrf/N158 ), .Q(
        \vrf/regTable[5][139] ) );
  LHQD1BWP \vrf/regTable_reg[5][140]  ( .E(n3584), .D(\vrf/N159 ), .Q(
        \vrf/regTable[5][140] ) );
  LHQD1BWP \vrf/regTable_reg[5][141]  ( .E(\vrf/N281 ), .D(\vrf/N160 ), .Q(
        \vrf/regTable[5][141] ) );
  LHQD1BWP \vrf/regTable_reg[5][142]  ( .E(n3584), .D(\vrf/N161 ), .Q(
        \vrf/regTable[5][142] ) );
  LHQD1BWP \vrf/regTable_reg[5][143]  ( .E(\vrf/N281 ), .D(\vrf/N162 ), .Q(
        \vrf/regTable[5][143] ) );
  LHQD1BWP \vrf/regTable_reg[5][144]  ( .E(n3584), .D(\vrf/N163 ), .Q(
        \vrf/regTable[5][144] ) );
  LHQD1BWP \vrf/regTable_reg[5][145]  ( .E(\vrf/N281 ), .D(\vrf/N164 ), .Q(
        \vrf/regTable[5][145] ) );
  LHQD1BWP \vrf/regTable_reg[5][146]  ( .E(n3584), .D(\vrf/N165 ), .Q(
        \vrf/regTable[5][146] ) );
  LHQD1BWP \vrf/regTable_reg[5][147]  ( .E(\vrf/N281 ), .D(\vrf/N166 ), .Q(
        \vrf/regTable[5][147] ) );
  LHQD1BWP \vrf/regTable_reg[5][148]  ( .E(n3584), .D(\vrf/N167 ), .Q(
        \vrf/regTable[5][148] ) );
  LHQD1BWP \vrf/regTable_reg[5][149]  ( .E(n3584), .D(\vrf/N168 ), .Q(
        \vrf/regTable[5][149] ) );
  LHQD1BWP \vrf/regTable_reg[5][150]  ( .E(n3584), .D(\vrf/N169 ), .Q(
        \vrf/regTable[5][150] ) );
  LHQD1BWP \vrf/regTable_reg[5][151]  ( .E(\vrf/N281 ), .D(\vrf/N170 ), .Q(
        \vrf/regTable[5][151] ) );
  LHQD1BWP \vrf/regTable_reg[5][152]  ( .E(n3584), .D(\vrf/N171 ), .Q(
        \vrf/regTable[5][152] ) );
  LHQD1BWP \vrf/regTable_reg[5][153]  ( .E(n3584), .D(\vrf/N172 ), .Q(
        \vrf/regTable[5][153] ) );
  LHQD1BWP \vrf/regTable_reg[5][154]  ( .E(n3584), .D(\vrf/N173 ), .Q(
        \vrf/regTable[5][154] ) );
  LHQD1BWP \vrf/regTable_reg[5][155]  ( .E(\vrf/N281 ), .D(\vrf/N174 ), .Q(
        \vrf/regTable[5][155] ) );
  LHQD1BWP \vrf/regTable_reg[5][156]  ( .E(n3584), .D(\vrf/N175 ), .Q(
        \vrf/regTable[5][156] ) );
  LHQD1BWP \vrf/regTable_reg[5][157]  ( .E(n3584), .D(\vrf/N176 ), .Q(
        \vrf/regTable[5][157] ) );
  LHQD1BWP \vrf/regTable_reg[5][158]  ( .E(n3584), .D(\vrf/N177 ), .Q(
        \vrf/regTable[5][158] ) );
  LHQD1BWP \vrf/regTable_reg[5][159]  ( .E(n3584), .D(\vrf/N178 ), .Q(
        \vrf/regTable[5][159] ) );
  LHQD1BWP \vrf/regTable_reg[5][160]  ( .E(\vrf/N281 ), .D(\vrf/N179 ), .Q(
        \vrf/regTable[5][160] ) );
  LHQD1BWP \vrf/regTable_reg[5][161]  ( .E(n3584), .D(\vrf/N180 ), .Q(
        \vrf/regTable[5][161] ) );
  LHQD1BWP \vrf/regTable_reg[5][162]  ( .E(n3584), .D(\vrf/N181 ), .Q(
        \vrf/regTable[5][162] ) );
  LHQD1BWP \vrf/regTable_reg[5][163]  ( .E(n3584), .D(\vrf/N182 ), .Q(
        \vrf/regTable[5][163] ) );
  LHQD1BWP \vrf/regTable_reg[5][164]  ( .E(\vrf/N281 ), .D(\vrf/N183 ), .Q(
        \vrf/regTable[5][164] ) );
  LHQD1BWP \vrf/regTable_reg[5][165]  ( .E(n3584), .D(\vrf/N184 ), .Q(
        \vrf/regTable[5][165] ) );
  LHQD1BWP \vrf/regTable_reg[5][166]  ( .E(n3584), .D(\vrf/N185 ), .Q(
        \vrf/regTable[5][166] ) );
  LHQD1BWP \vrf/regTable_reg[5][167]  ( .E(n3584), .D(\vrf/N186 ), .Q(
        \vrf/regTable[5][167] ) );
  LHQD1BWP \vrf/regTable_reg[5][168]  ( .E(\vrf/N281 ), .D(\vrf/N187 ), .Q(
        \vrf/regTable[5][168] ) );
  LHQD1BWP \vrf/regTable_reg[5][169]  ( .E(n3584), .D(\vrf/N188 ), .Q(
        \vrf/regTable[5][169] ) );
  LHQD1BWP \vrf/regTable_reg[5][170]  ( .E(n3584), .D(\vrf/N189 ), .Q(
        \vrf/regTable[5][170] ) );
  LHQD1BWP \vrf/regTable_reg[5][171]  ( .E(n3584), .D(\vrf/N190 ), .Q(
        \vrf/regTable[5][171] ) );
  LHQD1BWP \vrf/regTable_reg[5][172]  ( .E(n3584), .D(\vrf/N191 ), .Q(
        \vrf/regTable[5][172] ) );
  LHQD1BWP \vrf/regTable_reg[5][173]  ( .E(n3584), .D(\vrf/N192 ), .Q(
        \vrf/regTable[5][173] ) );
  LHQD1BWP \vrf/regTable_reg[5][174]  ( .E(\vrf/N281 ), .D(\vrf/N193 ), .Q(
        \vrf/regTable[5][174] ) );
  LHQD1BWP \vrf/regTable_reg[5][175]  ( .E(n3584), .D(\vrf/N194 ), .Q(
        \vrf/regTable[5][175] ) );
  LHQD1BWP \vrf/regTable_reg[5][176]  ( .E(n3584), .D(\vrf/N195 ), .Q(
        \vrf/regTable[5][176] ) );
  LHQD1BWP \vrf/regTable_reg[5][177]  ( .E(n3584), .D(\vrf/N196 ), .Q(
        \vrf/regTable[5][177] ) );
  LHQD1BWP \vrf/regTable_reg[5][178]  ( .E(n3584), .D(\vrf/N197 ), .Q(
        \vrf/regTable[5][178] ) );
  LHQD1BWP \vrf/regTable_reg[5][179]  ( .E(\vrf/N281 ), .D(\vrf/N198 ), .Q(
        \vrf/regTable[5][179] ) );
  LHQD1BWP \vrf/regTable_reg[5][180]  ( .E(n3584), .D(\vrf/N199 ), .Q(
        \vrf/regTable[5][180] ) );
  LHQD1BWP \vrf/regTable_reg[5][181]  ( .E(n3584), .D(\vrf/N200 ), .Q(
        \vrf/regTable[5][181] ) );
  LHQD1BWP \vrf/regTable_reg[5][182]  ( .E(n3584), .D(\vrf/N201 ), .Q(
        \vrf/regTable[5][182] ) );
  LHQD1BWP \vrf/regTable_reg[5][183]  ( .E(n3584), .D(\vrf/N202 ), .Q(
        \vrf/regTable[5][183] ) );
  LHQD1BWP \vrf/regTable_reg[5][184]  ( .E(n3584), .D(\vrf/N203 ), .Q(
        \vrf/regTable[5][184] ) );
  LHQD1BWP \vrf/regTable_reg[5][185]  ( .E(n3584), .D(\vrf/N204 ), .Q(
        \vrf/regTable[5][185] ) );
  LHQD1BWP \vrf/regTable_reg[5][186]  ( .E(n3584), .D(\vrf/N205 ), .Q(
        \vrf/regTable[5][186] ) );
  LHQD1BWP \vrf/regTable_reg[5][187]  ( .E(n3584), .D(\vrf/N206 ), .Q(
        \vrf/regTable[5][187] ) );
  LHQD1BWP \vrf/regTable_reg[5][188]  ( .E(n3584), .D(\vrf/N207 ), .Q(
        \vrf/regTable[5][188] ) );
  LHQD1BWP \vrf/regTable_reg[5][189]  ( .E(\vrf/N281 ), .D(\vrf/N208 ), .Q(
        \vrf/regTable[5][189] ) );
  LHQD1BWP \vrf/regTable_reg[5][190]  ( .E(n3584), .D(\vrf/N209 ), .Q(
        \vrf/regTable[5][190] ) );
  LHQD1BWP \vrf/regTable_reg[5][191]  ( .E(n3584), .D(\vrf/N210 ), .Q(
        \vrf/regTable[5][191] ) );
  LHQD1BWP \vrf/regTable_reg[5][192]  ( .E(n3584), .D(\vrf/N211 ), .Q(
        \vrf/regTable[5][192] ) );
  LHQD1BWP \vrf/regTable_reg[5][193]  ( .E(n3584), .D(\vrf/N212 ), .Q(
        \vrf/regTable[5][193] ) );
  LHQD1BWP \vrf/regTable_reg[5][194]  ( .E(\vrf/N281 ), .D(\vrf/N213 ), .Q(
        \vrf/regTable[5][194] ) );
  LHQD1BWP \vrf/regTable_reg[5][195]  ( .E(\vrf/N281 ), .D(\vrf/N214 ), .Q(
        \vrf/regTable[5][195] ) );
  LHQD1BWP \vrf/regTable_reg[5][196]  ( .E(n3584), .D(\vrf/N215 ), .Q(
        \vrf/regTable[5][196] ) );
  LHQD1BWP \vrf/regTable_reg[5][197]  ( .E(n3584), .D(\vrf/N216 ), .Q(
        \vrf/regTable[5][197] ) );
  LHQD1BWP \vrf/regTable_reg[5][198]  ( .E(n3584), .D(\vrf/N218 ), .Q(
        \vrf/regTable[5][198] ) );
  LHQD1BWP \vrf/regTable_reg[5][199]  ( .E(n3584), .D(\vrf/N219 ), .Q(
        \vrf/regTable[5][199] ) );
  LHQD1BWP \vrf/regTable_reg[5][200]  ( .E(n3584), .D(\vrf/N220 ), .Q(
        \vrf/regTable[5][200] ) );
  LHQD1BWP \vrf/regTable_reg[5][201]  ( .E(\vrf/N281 ), .D(\vrf/N221 ), .Q(
        \vrf/regTable[5][201] ) );
  LHQD1BWP \vrf/regTable_reg[5][202]  ( .E(n3584), .D(\vrf/N222 ), .Q(
        \vrf/regTable[5][202] ) );
  LHQD1BWP \vrf/regTable_reg[5][203]  ( .E(n3584), .D(\vrf/N223 ), .Q(
        \vrf/regTable[5][203] ) );
  LHQD1BWP \vrf/regTable_reg[5][204]  ( .E(\vrf/N281 ), .D(\vrf/N224 ), .Q(
        \vrf/regTable[5][204] ) );
  LHQD1BWP \vrf/regTable_reg[5][205]  ( .E(n3584), .D(\vrf/N225 ), .Q(
        \vrf/regTable[5][205] ) );
  LHQD1BWP \vrf/regTable_reg[5][206]  ( .E(\vrf/N281 ), .D(\vrf/N226 ), .Q(
        \vrf/regTable[5][206] ) );
  LHQD1BWP \vrf/regTable_reg[5][207]  ( .E(n3584), .D(\vrf/N227 ), .Q(
        \vrf/regTable[5][207] ) );
  LHQD1BWP \vrf/regTable_reg[5][208]  ( .E(n3584), .D(\vrf/N228 ), .Q(
        \vrf/regTable[5][208] ) );
  LHQD1BWP \vrf/regTable_reg[5][209]  ( .E(n3584), .D(\vrf/N229 ), .Q(
        \vrf/regTable[5][209] ) );
  LHQD1BWP \vrf/regTable_reg[5][210]  ( .E(n3584), .D(\vrf/N230 ), .Q(
        \vrf/regTable[5][210] ) );
  LHQD1BWP \vrf/regTable_reg[5][211]  ( .E(n3584), .D(\vrf/N231 ), .Q(
        \vrf/regTable[5][211] ) );
  LHQD1BWP \vrf/regTable_reg[5][212]  ( .E(n3584), .D(\vrf/N232 ), .Q(
        \vrf/regTable[5][212] ) );
  LHQD1BWP \vrf/regTable_reg[5][213]  ( .E(n3584), .D(\vrf/N233 ), .Q(
        \vrf/regTable[5][213] ) );
  LHQD1BWP \vrf/regTable_reg[5][214]  ( .E(n3584), .D(\vrf/N234 ), .Q(
        \vrf/regTable[5][214] ) );
  LHQD1BWP \vrf/regTable_reg[5][215]  ( .E(n3584), .D(\vrf/N235 ), .Q(
        \vrf/regTable[5][215] ) );
  LHQD1BWP \vrf/regTable_reg[5][216]  ( .E(n3584), .D(\vrf/N236 ), .Q(
        \vrf/regTable[5][216] ) );
  LHQD1BWP \vrf/regTable_reg[5][217]  ( .E(n3584), .D(\vrf/N237 ), .Q(
        \vrf/regTable[5][217] ) );
  LHQD1BWP \vrf/regTable_reg[5][218]  ( .E(n3584), .D(\vrf/N238 ), .Q(
        \vrf/regTable[5][218] ) );
  LHQD1BWP \vrf/regTable_reg[5][219]  ( .E(n3584), .D(\vrf/N239 ), .Q(
        \vrf/regTable[5][219] ) );
  LHQD1BWP \vrf/regTable_reg[5][220]  ( .E(n3584), .D(\vrf/N240 ), .Q(
        \vrf/regTable[5][220] ) );
  LHQD1BWP \vrf/regTable_reg[5][221]  ( .E(n3584), .D(\vrf/N241 ), .Q(
        \vrf/regTable[5][221] ) );
  LHQD1BWP \vrf/regTable_reg[5][222]  ( .E(n3584), .D(\vrf/N242 ), .Q(
        \vrf/regTable[5][222] ) );
  LHQD1BWP \vrf/regTable_reg[5][223]  ( .E(\vrf/N281 ), .D(\vrf/N243 ), .Q(
        \vrf/regTable[5][223] ) );
  LHQD1BWP \vrf/regTable_reg[5][224]  ( .E(n3584), .D(\vrf/N244 ), .Q(
        \vrf/regTable[5][224] ) );
  LHQD1BWP \vrf/regTable_reg[5][225]  ( .E(n3584), .D(\vrf/N245 ), .Q(
        \vrf/regTable[5][225] ) );
  LHQD1BWP \vrf/regTable_reg[5][226]  ( .E(n3584), .D(\vrf/N246 ), .Q(
        \vrf/regTable[5][226] ) );
  LHQD1BWP \vrf/regTable_reg[5][227]  ( .E(\vrf/N281 ), .D(\vrf/N247 ), .Q(
        \vrf/regTable[5][227] ) );
  LHQD1BWP \vrf/regTable_reg[5][228]  ( .E(n3584), .D(\vrf/N248 ), .Q(
        \vrf/regTable[5][228] ) );
  LHQD1BWP \vrf/regTable_reg[5][229]  ( .E(n3584), .D(\vrf/N249 ), .Q(
        \vrf/regTable[5][229] ) );
  LHQD1BWP \vrf/regTable_reg[5][230]  ( .E(n3584), .D(\vrf/N250 ), .Q(
        \vrf/regTable[5][230] ) );
  LHQD1BWP \vrf/regTable_reg[5][231]  ( .E(\vrf/N281 ), .D(\vrf/N251 ), .Q(
        \vrf/regTable[5][231] ) );
  LHQD1BWP \vrf/regTable_reg[5][232]  ( .E(n3584), .D(\vrf/N252 ), .Q(
        \vrf/regTable[5][232] ) );
  LHQD1BWP \vrf/regTable_reg[5][233]  ( .E(n3584), .D(\vrf/N253 ), .Q(
        \vrf/regTable[5][233] ) );
  LHQD1BWP \vrf/regTable_reg[5][234]  ( .E(n3584), .D(\vrf/N254 ), .Q(
        \vrf/regTable[5][234] ) );
  LHQD1BWP \vrf/regTable_reg[5][235]  ( .E(n3584), .D(\vrf/N255 ), .Q(
        \vrf/regTable[5][235] ) );
  LHQD1BWP \vrf/regTable_reg[5][236]  ( .E(n3584), .D(\vrf/N256 ), .Q(
        \vrf/regTable[5][236] ) );
  LHQD1BWP \vrf/regTable_reg[5][237]  ( .E(n3584), .D(\vrf/N257 ), .Q(
        \vrf/regTable[5][237] ) );
  LHQD1BWP \vrf/regTable_reg[5][238]  ( .E(n3584), .D(\vrf/N258 ), .Q(
        \vrf/regTable[5][238] ) );
  LHQD1BWP \vrf/regTable_reg[5][239]  ( .E(n3584), .D(\vrf/N259 ), .Q(
        \vrf/regTable[5][239] ) );
  LHQD1BWP \vrf/regTable_reg[5][240]  ( .E(n3584), .D(\vrf/N260 ), .Q(
        \vrf/regTable[5][240] ) );
  LHQD1BWP \vrf/regTable_reg[5][241]  ( .E(n3584), .D(\vrf/N261 ), .Q(
        \vrf/regTable[5][241] ) );
  LHQD1BWP \vrf/regTable_reg[5][242]  ( .E(n3584), .D(\vrf/N262 ), .Q(
        \vrf/regTable[5][242] ) );
  LHQD1BWP \vrf/regTable_reg[5][243]  ( .E(n3584), .D(\vrf/N263 ), .Q(
        \vrf/regTable[5][243] ) );
  LHQD1BWP \vrf/regTable_reg[5][244]  ( .E(n3584), .D(\vrf/N264 ), .Q(
        \vrf/regTable[5][244] ) );
  LHQD1BWP \vrf/regTable_reg[5][245]  ( .E(n3584), .D(\vrf/N265 ), .Q(
        \vrf/regTable[5][245] ) );
  LHQD1BWP \vrf/regTable_reg[5][246]  ( .E(n3584), .D(\vrf/N266 ), .Q(
        \vrf/regTable[5][246] ) );
  LHQD1BWP \vrf/regTable_reg[5][247]  ( .E(n3584), .D(\vrf/N267 ), .Q(
        \vrf/regTable[5][247] ) );
  LHQD1BWP \vrf/regTable_reg[5][248]  ( .E(n3584), .D(\vrf/N268 ), .Q(
        \vrf/regTable[5][248] ) );
  LHQD1BWP \vrf/regTable_reg[5][249]  ( .E(n3584), .D(\vrf/N269 ), .Q(
        \vrf/regTable[5][249] ) );
  LHQD1BWP \vrf/regTable_reg[5][250]  ( .E(n3584), .D(\vrf/N270 ), .Q(
        \vrf/regTable[5][250] ) );
  LHQD1BWP \vrf/regTable_reg[5][251]  ( .E(\vrf/N281 ), .D(\vrf/N271 ), .Q(
        \vrf/regTable[5][251] ) );
  LHQD1BWP \vrf/regTable_reg[5][252]  ( .E(n3584), .D(\vrf/N272 ), .Q(
        \vrf/regTable[5][252] ) );
  LHQD1BWP \vrf/regTable_reg[5][253]  ( .E(n3584), .D(\vrf/N273 ), .Q(
        \vrf/regTable[5][253] ) );
  LHQD1BWP \vrf/regTable_reg[5][254]  ( .E(n3584), .D(\vrf/N274 ), .Q(
        \vrf/regTable[5][254] ) );
  LHQD1BWP \vrf/regTable_reg[5][255]  ( .E(n3584), .D(\vrf/N275 ), .Q(
        \vrf/regTable[5][255] ) );
  LHQD1BWP \vrf/regTable_reg[4][0]  ( .E(n3586), .D(\vrf/N18 ), .Q(
        \vrf/regTable[4][0] ) );
  LHQD1BWP \vrf/regTable_reg[4][1]  ( .E(n3586), .D(\vrf/N19 ), .Q(
        \vrf/regTable[4][1] ) );
  LHQD1BWP \vrf/regTable_reg[4][2]  ( .E(n3586), .D(\vrf/N20 ), .Q(
        \vrf/regTable[4][2] ) );
  LHQD1BWP \vrf/regTable_reg[4][3]  ( .E(n3586), .D(\vrf/N21 ), .Q(
        \vrf/regTable[4][3] ) );
  LHQD1BWP \vrf/regTable_reg[4][4]  ( .E(n3586), .D(\vrf/N22 ), .Q(
        \vrf/regTable[4][4] ) );
  LHQD1BWP \vrf/regTable_reg[4][5]  ( .E(n3586), .D(\vrf/N23 ), .Q(
        \vrf/regTable[4][5] ) );
  LHQD1BWP \vrf/regTable_reg[4][6]  ( .E(n3586), .D(\vrf/N24 ), .Q(
        \vrf/regTable[4][6] ) );
  LHQD1BWP \vrf/regTable_reg[4][7]  ( .E(n3586), .D(\vrf/N25 ), .Q(
        \vrf/regTable[4][7] ) );
  LHQD1BWP \vrf/regTable_reg[4][8]  ( .E(n3586), .D(\vrf/N26 ), .Q(
        \vrf/regTable[4][8] ) );
  LHQD1BWP \vrf/regTable_reg[4][9]  ( .E(n3586), .D(\vrf/N27 ), .Q(
        \vrf/regTable[4][9] ) );
  LHQD1BWP \vrf/regTable_reg[4][10]  ( .E(n3586), .D(\vrf/N28 ), .Q(
        \vrf/regTable[4][10] ) );
  LHQD1BWP \vrf/regTable_reg[4][11]  ( .E(n3586), .D(\vrf/N29 ), .Q(
        \vrf/regTable[4][11] ) );
  LHQD1BWP \vrf/regTable_reg[4][12]  ( .E(n3586), .D(\vrf/N30 ), .Q(
        \vrf/regTable[4][12] ) );
  LHQD1BWP \vrf/regTable_reg[4][13]  ( .E(n3586), .D(\vrf/N31 ), .Q(
        \vrf/regTable[4][13] ) );
  LHQD1BWP \vrf/regTable_reg[4][14]  ( .E(n3586), .D(\vrf/N32 ), .Q(
        \vrf/regTable[4][14] ) );
  LHQD1BWP \vrf/regTable_reg[4][15]  ( .E(n3586), .D(\vrf/N33 ), .Q(
        \vrf/regTable[4][15] ) );
  LHQD1BWP \vrf/regTable_reg[4][16]  ( .E(n3586), .D(\vrf/N34 ), .Q(
        \vrf/regTable[4][16] ) );
  LHQD1BWP \vrf/regTable_reg[4][17]  ( .E(n3586), .D(\vrf/N35 ), .Q(
        \vrf/regTable[4][17] ) );
  LHQD1BWP \vrf/regTable_reg[4][18]  ( .E(n3586), .D(\vrf/N36 ), .Q(
        \vrf/regTable[4][18] ) );
  LHQD1BWP \vrf/regTable_reg[4][19]  ( .E(n3586), .D(\vrf/N37 ), .Q(
        \vrf/regTable[4][19] ) );
  LHQD1BWP \vrf/regTable_reg[4][20]  ( .E(n3586), .D(\vrf/N38 ), .Q(
        \vrf/regTable[4][20] ) );
  LHQD1BWP \vrf/regTable_reg[4][21]  ( .E(n3586), .D(\vrf/N39 ), .Q(
        \vrf/regTable[4][21] ) );
  LHQD1BWP \vrf/regTable_reg[4][22]  ( .E(n3586), .D(\vrf/N40 ), .Q(
        \vrf/regTable[4][22] ) );
  LHQD1BWP \vrf/regTable_reg[4][23]  ( .E(n3586), .D(\vrf/N41 ), .Q(
        \vrf/regTable[4][23] ) );
  LHQD1BWP \vrf/regTable_reg[4][24]  ( .E(n3586), .D(\vrf/N42 ), .Q(
        \vrf/regTable[4][24] ) );
  LHQD1BWP \vrf/regTable_reg[4][25]  ( .E(n3586), .D(\vrf/N43 ), .Q(
        \vrf/regTable[4][25] ) );
  LHQD1BWP \vrf/regTable_reg[4][26]  ( .E(n3586), .D(\vrf/N44 ), .Q(
        \vrf/regTable[4][26] ) );
  LHQD1BWP \vrf/regTable_reg[4][27]  ( .E(n3586), .D(\vrf/N45 ), .Q(
        \vrf/regTable[4][27] ) );
  LHQD1BWP \vrf/regTable_reg[4][28]  ( .E(n3586), .D(\vrf/N46 ), .Q(
        \vrf/regTable[4][28] ) );
  LHQD1BWP \vrf/regTable_reg[4][29]  ( .E(n3586), .D(\vrf/N47 ), .Q(
        \vrf/regTable[4][29] ) );
  LHQD1BWP \vrf/regTable_reg[4][30]  ( .E(n3586), .D(\vrf/N48 ), .Q(
        \vrf/regTable[4][30] ) );
  LHQD1BWP \vrf/regTable_reg[4][31]  ( .E(n3586), .D(\vrf/N49 ), .Q(
        \vrf/regTable[4][31] ) );
  LHQD1BWP \vrf/regTable_reg[4][32]  ( .E(n3586), .D(\vrf/N50 ), .Q(
        \vrf/regTable[4][32] ) );
  LHQD1BWP \vrf/regTable_reg[4][33]  ( .E(n3586), .D(\vrf/N51 ), .Q(
        \vrf/regTable[4][33] ) );
  LHQD1BWP \vrf/regTable_reg[4][34]  ( .E(n3586), .D(\vrf/N52 ), .Q(
        \vrf/regTable[4][34] ) );
  LHQD1BWP \vrf/regTable_reg[4][35]  ( .E(n3586), .D(\vrf/N53 ), .Q(
        \vrf/regTable[4][35] ) );
  LHQD1BWP \vrf/regTable_reg[4][36]  ( .E(n3586), .D(\vrf/N54 ), .Q(
        \vrf/regTable[4][36] ) );
  LHQD1BWP \vrf/regTable_reg[4][37]  ( .E(n3586), .D(\vrf/N55 ), .Q(
        \vrf/regTable[4][37] ) );
  LHQD1BWP \vrf/regTable_reg[4][38]  ( .E(n3586), .D(\vrf/N56 ), .Q(
        \vrf/regTable[4][38] ) );
  LHQD1BWP \vrf/regTable_reg[4][39]  ( .E(n3586), .D(\vrf/N57 ), .Q(
        \vrf/regTable[4][39] ) );
  LHQD1BWP \vrf/regTable_reg[4][40]  ( .E(n3586), .D(\vrf/N58 ), .Q(
        \vrf/regTable[4][40] ) );
  LHQD1BWP \vrf/regTable_reg[4][41]  ( .E(n3586), .D(\vrf/N59 ), .Q(
        \vrf/regTable[4][41] ) );
  LHQD1BWP \vrf/regTable_reg[4][42]  ( .E(n3586), .D(\vrf/N60 ), .Q(
        \vrf/regTable[4][42] ) );
  LHQD1BWP \vrf/regTable_reg[4][43]  ( .E(n3586), .D(\vrf/N61 ), .Q(
        \vrf/regTable[4][43] ) );
  LHQD1BWP \vrf/regTable_reg[4][44]  ( .E(n3586), .D(\vrf/N62 ), .Q(
        \vrf/regTable[4][44] ) );
  LHQD1BWP \vrf/regTable_reg[4][45]  ( .E(n3586), .D(\vrf/N63 ), .Q(
        \vrf/regTable[4][45] ) );
  LHQD1BWP \vrf/regTable_reg[4][46]  ( .E(n3586), .D(\vrf/N64 ), .Q(
        \vrf/regTable[4][46] ) );
  LHQD1BWP \vrf/regTable_reg[4][47]  ( .E(n3586), .D(\vrf/N65 ), .Q(
        \vrf/regTable[4][47] ) );
  LHQD1BWP \vrf/regTable_reg[4][48]  ( .E(n3586), .D(\vrf/N66 ), .Q(
        \vrf/regTable[4][48] ) );
  LHQD1BWP \vrf/regTable_reg[4][49]  ( .E(n3586), .D(\vrf/N67 ), .Q(
        \vrf/regTable[4][49] ) );
  LHQD1BWP \vrf/regTable_reg[4][50]  ( .E(n3586), .D(\vrf/N68 ), .Q(
        \vrf/regTable[4][50] ) );
  LHQD1BWP \vrf/regTable_reg[4][51]  ( .E(n3586), .D(\vrf/N69 ), .Q(
        \vrf/regTable[4][51] ) );
  LHQD1BWP \vrf/regTable_reg[4][52]  ( .E(n3586), .D(\vrf/N70 ), .Q(
        \vrf/regTable[4][52] ) );
  LHQD1BWP \vrf/regTable_reg[4][53]  ( .E(n3586), .D(\vrf/N71 ), .Q(
        \vrf/regTable[4][53] ) );
  LHQD1BWP \vrf/regTable_reg[4][54]  ( .E(n3586), .D(\vrf/N72 ), .Q(
        \vrf/regTable[4][54] ) );
  LHQD1BWP \vrf/regTable_reg[4][55]  ( .E(n3586), .D(\vrf/N73 ), .Q(
        \vrf/regTable[4][55] ) );
  LHQD1BWP \vrf/regTable_reg[4][56]  ( .E(n3586), .D(\vrf/N74 ), .Q(
        \vrf/regTable[4][56] ) );
  LHQD1BWP \vrf/regTable_reg[4][57]  ( .E(n3586), .D(\vrf/N75 ), .Q(
        \vrf/regTable[4][57] ) );
  LHQD1BWP \vrf/regTable_reg[4][58]  ( .E(n3586), .D(\vrf/N76 ), .Q(
        \vrf/regTable[4][58] ) );
  LHQD1BWP \vrf/regTable_reg[4][59]  ( .E(n3586), .D(\vrf/N77 ), .Q(
        \vrf/regTable[4][59] ) );
  LHQD1BWP \vrf/regTable_reg[4][60]  ( .E(n3586), .D(\vrf/N78 ), .Q(
        \vrf/regTable[4][60] ) );
  LHQD1BWP \vrf/regTable_reg[4][61]  ( .E(n3586), .D(\vrf/N79 ), .Q(
        \vrf/regTable[4][61] ) );
  LHQD1BWP \vrf/regTable_reg[4][62]  ( .E(n3586), .D(\vrf/N80 ), .Q(
        \vrf/regTable[4][62] ) );
  LHQD1BWP \vrf/regTable_reg[4][63]  ( .E(n3586), .D(\vrf/N81 ), .Q(
        \vrf/regTable[4][63] ) );
  LHQD1BWP \vrf/regTable_reg[4][64]  ( .E(n3586), .D(\vrf/N82 ), .Q(
        \vrf/regTable[4][64] ) );
  LHQD1BWP \vrf/regTable_reg[4][65]  ( .E(n3586), .D(\vrf/N83 ), .Q(
        \vrf/regTable[4][65] ) );
  LHQD1BWP \vrf/regTable_reg[4][66]  ( .E(n3586), .D(\vrf/N84 ), .Q(
        \vrf/regTable[4][66] ) );
  LHQD1BWP \vrf/regTable_reg[4][67]  ( .E(n3586), .D(\vrf/N85 ), .Q(
        \vrf/regTable[4][67] ) );
  LHQD1BWP \vrf/regTable_reg[4][68]  ( .E(n3586), .D(\vrf/N86 ), .Q(
        \vrf/regTable[4][68] ) );
  LHQD1BWP \vrf/regTable_reg[4][69]  ( .E(n3586), .D(\vrf/N87 ), .Q(
        \vrf/regTable[4][69] ) );
  LHQD1BWP \vrf/regTable_reg[4][70]  ( .E(n3586), .D(\vrf/N88 ), .Q(
        \vrf/regTable[4][70] ) );
  LHQD1BWP \vrf/regTable_reg[4][71]  ( .E(n3586), .D(\vrf/N89 ), .Q(
        \vrf/regTable[4][71] ) );
  LHQD1BWP \vrf/regTable_reg[4][72]  ( .E(n3586), .D(\vrf/N90 ), .Q(
        \vrf/regTable[4][72] ) );
  LHQD1BWP \vrf/regTable_reg[4][73]  ( .E(n3586), .D(\vrf/N91 ), .Q(
        \vrf/regTable[4][73] ) );
  LHQD1BWP \vrf/regTable_reg[4][74]  ( .E(n3586), .D(\vrf/N92 ), .Q(
        \vrf/regTable[4][74] ) );
  LHQD1BWP \vrf/regTable_reg[4][75]  ( .E(n3586), .D(\vrf/N93 ), .Q(
        \vrf/regTable[4][75] ) );
  LHQD1BWP \vrf/regTable_reg[4][76]  ( .E(n3586), .D(\vrf/N94 ), .Q(
        \vrf/regTable[4][76] ) );
  LHQD1BWP \vrf/regTable_reg[4][77]  ( .E(n3586), .D(\vrf/N95 ), .Q(
        \vrf/regTable[4][77] ) );
  LHQD1BWP \vrf/regTable_reg[4][78]  ( .E(n3586), .D(\vrf/N96 ), .Q(
        \vrf/regTable[4][78] ) );
  LHQD1BWP \vrf/regTable_reg[4][79]  ( .E(n3586), .D(\vrf/N97 ), .Q(
        \vrf/regTable[4][79] ) );
  LHQD1BWP \vrf/regTable_reg[4][80]  ( .E(n3586), .D(\vrf/N98 ), .Q(
        \vrf/regTable[4][80] ) );
  LHQD1BWP \vrf/regTable_reg[4][81]  ( .E(n3586), .D(\vrf/N99 ), .Q(
        \vrf/regTable[4][81] ) );
  LHQD1BWP \vrf/regTable_reg[4][82]  ( .E(n3586), .D(\vrf/N100 ), .Q(
        \vrf/regTable[4][82] ) );
  LHQD1BWP \vrf/regTable_reg[4][83]  ( .E(n3586), .D(\vrf/N101 ), .Q(
        \vrf/regTable[4][83] ) );
  LHQD1BWP \vrf/regTable_reg[4][84]  ( .E(n3586), .D(\vrf/N102 ), .Q(
        \vrf/regTable[4][84] ) );
  LHQD1BWP \vrf/regTable_reg[4][85]  ( .E(n3586), .D(\vrf/N103 ), .Q(
        \vrf/regTable[4][85] ) );
  LHQD1BWP \vrf/regTable_reg[4][86]  ( .E(n3586), .D(\vrf/N104 ), .Q(
        \vrf/regTable[4][86] ) );
  LHQD1BWP \vrf/regTable_reg[4][87]  ( .E(n3586), .D(\vrf/N105 ), .Q(
        \vrf/regTable[4][87] ) );
  LHQD1BWP \vrf/regTable_reg[4][88]  ( .E(n3586), .D(\vrf/N106 ), .Q(
        \vrf/regTable[4][88] ) );
  LHQD1BWP \vrf/regTable_reg[4][89]  ( .E(n3586), .D(\vrf/N107 ), .Q(
        \vrf/regTable[4][89] ) );
  LHQD1BWP \vrf/regTable_reg[4][90]  ( .E(n3586), .D(\vrf/N108 ), .Q(
        \vrf/regTable[4][90] ) );
  LHQD1BWP \vrf/regTable_reg[4][91]  ( .E(n3586), .D(\vrf/N109 ), .Q(
        \vrf/regTable[4][91] ) );
  LHQD1BWP \vrf/regTable_reg[4][92]  ( .E(n3586), .D(\vrf/N110 ), .Q(
        \vrf/regTable[4][92] ) );
  LHQD1BWP \vrf/regTable_reg[4][93]  ( .E(n3586), .D(\vrf/N111 ), .Q(
        \vrf/regTable[4][93] ) );
  LHQD1BWP \vrf/regTable_reg[4][94]  ( .E(n3586), .D(\vrf/N112 ), .Q(
        \vrf/regTable[4][94] ) );
  LHQD1BWP \vrf/regTable_reg[4][95]  ( .E(n3586), .D(\vrf/N113 ), .Q(
        \vrf/regTable[4][95] ) );
  LHQD1BWP \vrf/regTable_reg[4][96]  ( .E(n3586), .D(\vrf/N114 ), .Q(
        \vrf/regTable[4][96] ) );
  LHQD1BWP \vrf/regTable_reg[4][97]  ( .E(n3586), .D(\vrf/N115 ), .Q(
        \vrf/regTable[4][97] ) );
  LHQD1BWP \vrf/regTable_reg[4][98]  ( .E(n3586), .D(\vrf/N116 ), .Q(
        \vrf/regTable[4][98] ) );
  LHQD1BWP \vrf/regTable_reg[4][99]  ( .E(n3586), .D(\vrf/N118 ), .Q(
        \vrf/regTable[4][99] ) );
  LHQD1BWP \vrf/regTable_reg[4][100]  ( .E(n3586), .D(\vrf/N119 ), .Q(
        \vrf/regTable[4][100] ) );
  LHQD1BWP \vrf/regTable_reg[4][101]  ( .E(n3586), .D(\vrf/N120 ), .Q(
        \vrf/regTable[4][101] ) );
  LHQD1BWP \vrf/regTable_reg[4][102]  ( .E(n3586), .D(\vrf/N121 ), .Q(
        \vrf/regTable[4][102] ) );
  LHQD1BWP \vrf/regTable_reg[4][103]  ( .E(n3586), .D(\vrf/N122 ), .Q(
        \vrf/regTable[4][103] ) );
  LHQD1BWP \vrf/regTable_reg[4][104]  ( .E(n3586), .D(\vrf/N123 ), .Q(
        \vrf/regTable[4][104] ) );
  LHQD1BWP \vrf/regTable_reg[4][105]  ( .E(n3586), .D(\vrf/N124 ), .Q(
        \vrf/regTable[4][105] ) );
  LHQD1BWP \vrf/regTable_reg[4][106]  ( .E(n3586), .D(\vrf/N125 ), .Q(
        \vrf/regTable[4][106] ) );
  LHQD1BWP \vrf/regTable_reg[4][107]  ( .E(n3586), .D(\vrf/N126 ), .Q(
        \vrf/regTable[4][107] ) );
  LHQD1BWP \vrf/regTable_reg[4][108]  ( .E(n3586), .D(\vrf/N127 ), .Q(
        \vrf/regTable[4][108] ) );
  LHQD1BWP \vrf/regTable_reg[4][109]  ( .E(n3586), .D(\vrf/N128 ), .Q(
        \vrf/regTable[4][109] ) );
  LHQD1BWP \vrf/regTable_reg[4][110]  ( .E(n3586), .D(\vrf/N129 ), .Q(
        \vrf/regTable[4][110] ) );
  LHQD1BWP \vrf/regTable_reg[4][111]  ( .E(n3586), .D(\vrf/N130 ), .Q(
        \vrf/regTable[4][111] ) );
  LHQD1BWP \vrf/regTable_reg[4][112]  ( .E(n3586), .D(\vrf/N131 ), .Q(
        \vrf/regTable[4][112] ) );
  LHQD1BWP \vrf/regTable_reg[4][113]  ( .E(n3586), .D(\vrf/N132 ), .Q(
        \vrf/regTable[4][113] ) );
  LHQD1BWP \vrf/regTable_reg[4][114]  ( .E(n3586), .D(\vrf/N133 ), .Q(
        \vrf/regTable[4][114] ) );
  LHQD1BWP \vrf/regTable_reg[4][115]  ( .E(n3586), .D(\vrf/N134 ), .Q(
        \vrf/regTable[4][115] ) );
  LHQD1BWP \vrf/regTable_reg[4][116]  ( .E(n3586), .D(\vrf/N135 ), .Q(
        \vrf/regTable[4][116] ) );
  LHQD1BWP \vrf/regTable_reg[4][117]  ( .E(n3586), .D(\vrf/N136 ), .Q(
        \vrf/regTable[4][117] ) );
  LHQD1BWP \vrf/regTable_reg[4][118]  ( .E(n3586), .D(\vrf/N137 ), .Q(
        \vrf/regTable[4][118] ) );
  LHQD1BWP \vrf/regTable_reg[4][119]  ( .E(n3586), .D(\vrf/N138 ), .Q(
        \vrf/regTable[4][119] ) );
  LHQD1BWP \vrf/regTable_reg[4][120]  ( .E(n3586), .D(\vrf/N139 ), .Q(
        \vrf/regTable[4][120] ) );
  LHQD1BWP \vrf/regTable_reg[4][121]  ( .E(n3586), .D(\vrf/N140 ), .Q(
        \vrf/regTable[4][121] ) );
  LHQD1BWP \vrf/regTable_reg[4][122]  ( .E(n3586), .D(\vrf/N141 ), .Q(
        \vrf/regTable[4][122] ) );
  LHQD1BWP \vrf/regTable_reg[4][123]  ( .E(n3586), .D(\vrf/N142 ), .Q(
        \vrf/regTable[4][123] ) );
  LHQD1BWP \vrf/regTable_reg[4][124]  ( .E(n3586), .D(\vrf/N143 ), .Q(
        \vrf/regTable[4][124] ) );
  LHQD1BWP \vrf/regTable_reg[4][125]  ( .E(n3586), .D(\vrf/N144 ), .Q(
        \vrf/regTable[4][125] ) );
  LHQD1BWP \vrf/regTable_reg[4][126]  ( .E(n3586), .D(\vrf/N145 ), .Q(
        \vrf/regTable[4][126] ) );
  LHQD1BWP \vrf/regTable_reg[4][127]  ( .E(n3586), .D(\vrf/N146 ), .Q(
        \vrf/regTable[4][127] ) );
  LHQD1BWP \vrf/regTable_reg[4][128]  ( .E(n3586), .D(\vrf/N147 ), .Q(
        \vrf/regTable[4][128] ) );
  LHQD1BWP \vrf/regTable_reg[4][129]  ( .E(n3586), .D(\vrf/N148 ), .Q(
        \vrf/regTable[4][129] ) );
  LHQD1BWP \vrf/regTable_reg[4][130]  ( .E(n3586), .D(\vrf/N149 ), .Q(
        \vrf/regTable[4][130] ) );
  LHQD1BWP \vrf/regTable_reg[4][131]  ( .E(n3586), .D(\vrf/N150 ), .Q(
        \vrf/regTable[4][131] ) );
  LHQD1BWP \vrf/regTable_reg[4][132]  ( .E(n3586), .D(\vrf/N151 ), .Q(
        \vrf/regTable[4][132] ) );
  LHQD1BWP \vrf/regTable_reg[4][133]  ( .E(n3586), .D(\vrf/N152 ), .Q(
        \vrf/regTable[4][133] ) );
  LHQD1BWP \vrf/regTable_reg[4][134]  ( .E(n3586), .D(\vrf/N153 ), .Q(
        \vrf/regTable[4][134] ) );
  LHQD1BWP \vrf/regTable_reg[4][135]  ( .E(n3586), .D(\vrf/N154 ), .Q(
        \vrf/regTable[4][135] ) );
  LHQD1BWP \vrf/regTable_reg[4][136]  ( .E(n3586), .D(\vrf/N155 ), .Q(
        \vrf/regTable[4][136] ) );
  LHQD1BWP \vrf/regTable_reg[4][137]  ( .E(\vrf/N284 ), .D(\vrf/N156 ), .Q(
        \vrf/regTable[4][137] ) );
  LHQD1BWP \vrf/regTable_reg[4][138]  ( .E(n3586), .D(\vrf/N157 ), .Q(
        \vrf/regTable[4][138] ) );
  LHQD1BWP \vrf/regTable_reg[4][139]  ( .E(\vrf/N284 ), .D(\vrf/N158 ), .Q(
        \vrf/regTable[4][139] ) );
  LHQD1BWP \vrf/regTable_reg[4][140]  ( .E(n3586), .D(\vrf/N159 ), .Q(
        \vrf/regTable[4][140] ) );
  LHQD1BWP \vrf/regTable_reg[4][141]  ( .E(\vrf/N284 ), .D(\vrf/N160 ), .Q(
        \vrf/regTable[4][141] ) );
  LHQD1BWP \vrf/regTable_reg[4][142]  ( .E(n3586), .D(\vrf/N161 ), .Q(
        \vrf/regTable[4][142] ) );
  LHQD1BWP \vrf/regTable_reg[4][143]  ( .E(\vrf/N284 ), .D(\vrf/N162 ), .Q(
        \vrf/regTable[4][143] ) );
  LHQD1BWP \vrf/regTable_reg[4][144]  ( .E(n3586), .D(\vrf/N163 ), .Q(
        \vrf/regTable[4][144] ) );
  LHQD1BWP \vrf/regTable_reg[4][145]  ( .E(\vrf/N284 ), .D(\vrf/N164 ), .Q(
        \vrf/regTable[4][145] ) );
  LHQD1BWP \vrf/regTable_reg[4][146]  ( .E(n3586), .D(\vrf/N165 ), .Q(
        \vrf/regTable[4][146] ) );
  LHQD1BWP \vrf/regTable_reg[4][147]  ( .E(\vrf/N284 ), .D(\vrf/N166 ), .Q(
        \vrf/regTable[4][147] ) );
  LHQD1BWP \vrf/regTable_reg[4][148]  ( .E(n3586), .D(\vrf/N167 ), .Q(
        \vrf/regTable[4][148] ) );
  LHQD1BWP \vrf/regTable_reg[4][149]  ( .E(n3586), .D(\vrf/N168 ), .Q(
        \vrf/regTable[4][149] ) );
  LHQD1BWP \vrf/regTable_reg[4][150]  ( .E(n3586), .D(\vrf/N169 ), .Q(
        \vrf/regTable[4][150] ) );
  LHQD1BWP \vrf/regTable_reg[4][151]  ( .E(\vrf/N284 ), .D(\vrf/N170 ), .Q(
        \vrf/regTable[4][151] ) );
  LHQD1BWP \vrf/regTable_reg[4][152]  ( .E(n3586), .D(\vrf/N171 ), .Q(
        \vrf/regTable[4][152] ) );
  LHQD1BWP \vrf/regTable_reg[4][153]  ( .E(n3586), .D(\vrf/N172 ), .Q(
        \vrf/regTable[4][153] ) );
  LHQD1BWP \vrf/regTable_reg[4][154]  ( .E(n3586), .D(\vrf/N173 ), .Q(
        \vrf/regTable[4][154] ) );
  LHQD1BWP \vrf/regTable_reg[4][155]  ( .E(\vrf/N284 ), .D(\vrf/N174 ), .Q(
        \vrf/regTable[4][155] ) );
  LHQD1BWP \vrf/regTable_reg[4][156]  ( .E(n3586), .D(\vrf/N175 ), .Q(
        \vrf/regTable[4][156] ) );
  LHQD1BWP \vrf/regTable_reg[4][157]  ( .E(n3586), .D(\vrf/N176 ), .Q(
        \vrf/regTable[4][157] ) );
  LHQD1BWP \vrf/regTable_reg[4][158]  ( .E(n3586), .D(\vrf/N177 ), .Q(
        \vrf/regTable[4][158] ) );
  LHQD1BWP \vrf/regTable_reg[4][159]  ( .E(n3586), .D(\vrf/N178 ), .Q(
        \vrf/regTable[4][159] ) );
  LHQD1BWP \vrf/regTable_reg[4][160]  ( .E(\vrf/N284 ), .D(\vrf/N179 ), .Q(
        \vrf/regTable[4][160] ) );
  LHQD1BWP \vrf/regTable_reg[4][161]  ( .E(n3586), .D(\vrf/N180 ), .Q(
        \vrf/regTable[4][161] ) );
  LHQD1BWP \vrf/regTable_reg[4][162]  ( .E(n3586), .D(\vrf/N181 ), .Q(
        \vrf/regTable[4][162] ) );
  LHQD1BWP \vrf/regTable_reg[4][163]  ( .E(n3586), .D(\vrf/N182 ), .Q(
        \vrf/regTable[4][163] ) );
  LHQD1BWP \vrf/regTable_reg[4][164]  ( .E(\vrf/N284 ), .D(\vrf/N183 ), .Q(
        \vrf/regTable[4][164] ) );
  LHQD1BWP \vrf/regTable_reg[4][165]  ( .E(n3586), .D(\vrf/N184 ), .Q(
        \vrf/regTable[4][165] ) );
  LHQD1BWP \vrf/regTable_reg[4][166]  ( .E(n3586), .D(\vrf/N185 ), .Q(
        \vrf/regTable[4][166] ) );
  LHQD1BWP \vrf/regTable_reg[4][167]  ( .E(n3586), .D(\vrf/N186 ), .Q(
        \vrf/regTable[4][167] ) );
  LHQD1BWP \vrf/regTable_reg[4][168]  ( .E(\vrf/N284 ), .D(\vrf/N187 ), .Q(
        \vrf/regTable[4][168] ) );
  LHQD1BWP \vrf/regTable_reg[4][169]  ( .E(n3586), .D(\vrf/N188 ), .Q(
        \vrf/regTable[4][169] ) );
  LHQD1BWP \vrf/regTable_reg[4][170]  ( .E(n3586), .D(\vrf/N189 ), .Q(
        \vrf/regTable[4][170] ) );
  LHQD1BWP \vrf/regTable_reg[4][171]  ( .E(n3586), .D(\vrf/N190 ), .Q(
        \vrf/regTable[4][171] ) );
  LHQD1BWP \vrf/regTable_reg[4][172]  ( .E(n3586), .D(\vrf/N191 ), .Q(
        \vrf/regTable[4][172] ) );
  LHQD1BWP \vrf/regTable_reg[4][173]  ( .E(n3586), .D(\vrf/N192 ), .Q(
        \vrf/regTable[4][173] ) );
  LHQD1BWP \vrf/regTable_reg[4][174]  ( .E(\vrf/N284 ), .D(\vrf/N193 ), .Q(
        \vrf/regTable[4][174] ) );
  LHQD1BWP \vrf/regTable_reg[4][175]  ( .E(n3586), .D(\vrf/N194 ), .Q(
        \vrf/regTable[4][175] ) );
  LHQD1BWP \vrf/regTable_reg[4][176]  ( .E(n3586), .D(\vrf/N195 ), .Q(
        \vrf/regTable[4][176] ) );
  LHQD1BWP \vrf/regTable_reg[4][177]  ( .E(n3586), .D(\vrf/N196 ), .Q(
        \vrf/regTable[4][177] ) );
  LHQD1BWP \vrf/regTable_reg[4][178]  ( .E(n3586), .D(\vrf/N197 ), .Q(
        \vrf/regTable[4][178] ) );
  LHQD1BWP \vrf/regTable_reg[4][179]  ( .E(\vrf/N284 ), .D(\vrf/N198 ), .Q(
        \vrf/regTable[4][179] ) );
  LHQD1BWP \vrf/regTable_reg[4][180]  ( .E(n3586), .D(\vrf/N199 ), .Q(
        \vrf/regTable[4][180] ) );
  LHQD1BWP \vrf/regTable_reg[4][181]  ( .E(n3586), .D(\vrf/N200 ), .Q(
        \vrf/regTable[4][181] ) );
  LHQD1BWP \vrf/regTable_reg[4][182]  ( .E(n3586), .D(\vrf/N201 ), .Q(
        \vrf/regTable[4][182] ) );
  LHQD1BWP \vrf/regTable_reg[4][183]  ( .E(n3586), .D(\vrf/N202 ), .Q(
        \vrf/regTable[4][183] ) );
  LHQD1BWP \vrf/regTable_reg[4][184]  ( .E(n3586), .D(\vrf/N203 ), .Q(
        \vrf/regTable[4][184] ) );
  LHQD1BWP \vrf/regTable_reg[4][185]  ( .E(n3586), .D(\vrf/N204 ), .Q(
        \vrf/regTable[4][185] ) );
  LHQD1BWP \vrf/regTable_reg[4][186]  ( .E(n3586), .D(\vrf/N205 ), .Q(
        \vrf/regTable[4][186] ) );
  LHQD1BWP \vrf/regTable_reg[4][187]  ( .E(n3586), .D(\vrf/N206 ), .Q(
        \vrf/regTable[4][187] ) );
  LHQD1BWP \vrf/regTable_reg[4][188]  ( .E(n3586), .D(\vrf/N207 ), .Q(
        \vrf/regTable[4][188] ) );
  LHQD1BWP \vrf/regTable_reg[4][189]  ( .E(\vrf/N284 ), .D(\vrf/N208 ), .Q(
        \vrf/regTable[4][189] ) );
  LHQD1BWP \vrf/regTable_reg[4][190]  ( .E(n3586), .D(\vrf/N209 ), .Q(
        \vrf/regTable[4][190] ) );
  LHQD1BWP \vrf/regTable_reg[4][191]  ( .E(n3586), .D(\vrf/N210 ), .Q(
        \vrf/regTable[4][191] ) );
  LHQD1BWP \vrf/regTable_reg[4][192]  ( .E(n3586), .D(\vrf/N211 ), .Q(
        \vrf/regTable[4][192] ) );
  LHQD1BWP \vrf/regTable_reg[4][193]  ( .E(n3586), .D(\vrf/N212 ), .Q(
        \vrf/regTable[4][193] ) );
  LHQD1BWP \vrf/regTable_reg[4][194]  ( .E(\vrf/N284 ), .D(\vrf/N213 ), .Q(
        \vrf/regTable[4][194] ) );
  LHQD1BWP \vrf/regTable_reg[4][195]  ( .E(\vrf/N284 ), .D(\vrf/N214 ), .Q(
        \vrf/regTable[4][195] ) );
  LHQD1BWP \vrf/regTable_reg[4][196]  ( .E(n3586), .D(\vrf/N215 ), .Q(
        \vrf/regTable[4][196] ) );
  LHQD1BWP \vrf/regTable_reg[4][197]  ( .E(n3586), .D(\vrf/N216 ), .Q(
        \vrf/regTable[4][197] ) );
  LHQD1BWP \vrf/regTable_reg[4][198]  ( .E(n3586), .D(\vrf/N218 ), .Q(
        \vrf/regTable[4][198] ) );
  LHQD1BWP \vrf/regTable_reg[4][199]  ( .E(n3586), .D(\vrf/N219 ), .Q(
        \vrf/regTable[4][199] ) );
  LHQD1BWP \vrf/regTable_reg[4][200]  ( .E(n3586), .D(\vrf/N220 ), .Q(
        \vrf/regTable[4][200] ) );
  LHQD1BWP \vrf/regTable_reg[4][201]  ( .E(\vrf/N284 ), .D(\vrf/N221 ), .Q(
        \vrf/regTable[4][201] ) );
  LHQD1BWP \vrf/regTable_reg[4][202]  ( .E(n3586), .D(\vrf/N222 ), .Q(
        \vrf/regTable[4][202] ) );
  LHQD1BWP \vrf/regTable_reg[4][203]  ( .E(n3586), .D(\vrf/N223 ), .Q(
        \vrf/regTable[4][203] ) );
  LHQD1BWP \vrf/regTable_reg[4][204]  ( .E(\vrf/N284 ), .D(\vrf/N224 ), .Q(
        \vrf/regTable[4][204] ) );
  LHQD1BWP \vrf/regTable_reg[4][205]  ( .E(n3586), .D(\vrf/N225 ), .Q(
        \vrf/regTable[4][205] ) );
  LHQD1BWP \vrf/regTable_reg[4][206]  ( .E(\vrf/N284 ), .D(\vrf/N226 ), .Q(
        \vrf/regTable[4][206] ) );
  LHQD1BWP \vrf/regTable_reg[4][207]  ( .E(n3586), .D(\vrf/N227 ), .Q(
        \vrf/regTable[4][207] ) );
  LHQD1BWP \vrf/regTable_reg[4][208]  ( .E(n3586), .D(\vrf/N228 ), .Q(
        \vrf/regTable[4][208] ) );
  LHQD1BWP \vrf/regTable_reg[4][209]  ( .E(n3586), .D(\vrf/N229 ), .Q(
        \vrf/regTable[4][209] ) );
  LHQD1BWP \vrf/regTable_reg[4][210]  ( .E(n3586), .D(\vrf/N230 ), .Q(
        \vrf/regTable[4][210] ) );
  LHQD1BWP \vrf/regTable_reg[4][211]  ( .E(n3586), .D(\vrf/N231 ), .Q(
        \vrf/regTable[4][211] ) );
  LHQD1BWP \vrf/regTable_reg[4][212]  ( .E(n3586), .D(\vrf/N232 ), .Q(
        \vrf/regTable[4][212] ) );
  LHQD1BWP \vrf/regTable_reg[4][213]  ( .E(n3586), .D(\vrf/N233 ), .Q(
        \vrf/regTable[4][213] ) );
  LHQD1BWP \vrf/regTable_reg[4][214]  ( .E(n3586), .D(\vrf/N234 ), .Q(
        \vrf/regTable[4][214] ) );
  LHQD1BWP \vrf/regTable_reg[4][215]  ( .E(n3586), .D(\vrf/N235 ), .Q(
        \vrf/regTable[4][215] ) );
  LHQD1BWP \vrf/regTable_reg[4][216]  ( .E(n3586), .D(\vrf/N236 ), .Q(
        \vrf/regTable[4][216] ) );
  LHQD1BWP \vrf/regTable_reg[4][217]  ( .E(n3586), .D(\vrf/N237 ), .Q(
        \vrf/regTable[4][217] ) );
  LHQD1BWP \vrf/regTable_reg[4][218]  ( .E(n3586), .D(\vrf/N238 ), .Q(
        \vrf/regTable[4][218] ) );
  LHQD1BWP \vrf/regTable_reg[4][219]  ( .E(n3586), .D(\vrf/N239 ), .Q(
        \vrf/regTable[4][219] ) );
  LHQD1BWP \vrf/regTable_reg[4][220]  ( .E(n3586), .D(\vrf/N240 ), .Q(
        \vrf/regTable[4][220] ) );
  LHQD1BWP \vrf/regTable_reg[4][221]  ( .E(n3586), .D(\vrf/N241 ), .Q(
        \vrf/regTable[4][221] ) );
  LHQD1BWP \vrf/regTable_reg[4][222]  ( .E(n3586), .D(\vrf/N242 ), .Q(
        \vrf/regTable[4][222] ) );
  LHQD1BWP \vrf/regTable_reg[4][223]  ( .E(\vrf/N284 ), .D(\vrf/N243 ), .Q(
        \vrf/regTable[4][223] ) );
  LHQD1BWP \vrf/regTable_reg[4][224]  ( .E(n3586), .D(\vrf/N244 ), .Q(
        \vrf/regTable[4][224] ) );
  LHQD1BWP \vrf/regTable_reg[4][225]  ( .E(n3586), .D(\vrf/N245 ), .Q(
        \vrf/regTable[4][225] ) );
  LHQD1BWP \vrf/regTable_reg[4][226]  ( .E(n3586), .D(\vrf/N246 ), .Q(
        \vrf/regTable[4][226] ) );
  LHQD1BWP \vrf/regTable_reg[4][227]  ( .E(\vrf/N284 ), .D(\vrf/N247 ), .Q(
        \vrf/regTable[4][227] ) );
  LHQD1BWP \vrf/regTable_reg[4][228]  ( .E(n3586), .D(\vrf/N248 ), .Q(
        \vrf/regTable[4][228] ) );
  LHQD1BWP \vrf/regTable_reg[4][229]  ( .E(n3586), .D(\vrf/N249 ), .Q(
        \vrf/regTable[4][229] ) );
  LHQD1BWP \vrf/regTable_reg[4][230]  ( .E(n3586), .D(\vrf/N250 ), .Q(
        \vrf/regTable[4][230] ) );
  LHQD1BWP \vrf/regTable_reg[4][231]  ( .E(\vrf/N284 ), .D(\vrf/N251 ), .Q(
        \vrf/regTable[4][231] ) );
  LHQD1BWP \vrf/regTable_reg[4][232]  ( .E(n3586), .D(\vrf/N252 ), .Q(
        \vrf/regTable[4][232] ) );
  LHQD1BWP \vrf/regTable_reg[4][233]  ( .E(n3586), .D(\vrf/N253 ), .Q(
        \vrf/regTable[4][233] ) );
  LHQD1BWP \vrf/regTable_reg[4][234]  ( .E(n3586), .D(\vrf/N254 ), .Q(
        \vrf/regTable[4][234] ) );
  LHQD1BWP \vrf/regTable_reg[4][235]  ( .E(n3586), .D(\vrf/N255 ), .Q(
        \vrf/regTable[4][235] ) );
  LHQD1BWP \vrf/regTable_reg[4][236]  ( .E(n3586), .D(\vrf/N256 ), .Q(
        \vrf/regTable[4][236] ) );
  LHQD1BWP \vrf/regTable_reg[4][237]  ( .E(n3586), .D(\vrf/N257 ), .Q(
        \vrf/regTable[4][237] ) );
  LHQD1BWP \vrf/regTable_reg[4][238]  ( .E(n3586), .D(\vrf/N258 ), .Q(
        \vrf/regTable[4][238] ) );
  LHQD1BWP \vrf/regTable_reg[4][239]  ( .E(n3586), .D(\vrf/N259 ), .Q(
        \vrf/regTable[4][239] ) );
  LHQD1BWP \vrf/regTable_reg[4][240]  ( .E(n3586), .D(\vrf/N260 ), .Q(
        \vrf/regTable[4][240] ) );
  LHQD1BWP \vrf/regTable_reg[4][241]  ( .E(n3586), .D(\vrf/N261 ), .Q(
        \vrf/regTable[4][241] ) );
  LHQD1BWP \vrf/regTable_reg[4][242]  ( .E(n3586), .D(\vrf/N262 ), .Q(
        \vrf/regTable[4][242] ) );
  LHQD1BWP \vrf/regTable_reg[4][243]  ( .E(n3586), .D(\vrf/N263 ), .Q(
        \vrf/regTable[4][243] ) );
  LHQD1BWP \vrf/regTable_reg[4][244]  ( .E(n3586), .D(\vrf/N264 ), .Q(
        \vrf/regTable[4][244] ) );
  LHQD1BWP \vrf/regTable_reg[4][245]  ( .E(n3586), .D(\vrf/N265 ), .Q(
        \vrf/regTable[4][245] ) );
  LHQD1BWP \vrf/regTable_reg[4][246]  ( .E(n3586), .D(\vrf/N266 ), .Q(
        \vrf/regTable[4][246] ) );
  LHQD1BWP \vrf/regTable_reg[4][247]  ( .E(n3586), .D(\vrf/N267 ), .Q(
        \vrf/regTable[4][247] ) );
  LHQD1BWP \vrf/regTable_reg[4][248]  ( .E(n3586), .D(\vrf/N268 ), .Q(
        \vrf/regTable[4][248] ) );
  LHQD1BWP \vrf/regTable_reg[4][249]  ( .E(n3586), .D(\vrf/N269 ), .Q(
        \vrf/regTable[4][249] ) );
  LHQD1BWP \vrf/regTable_reg[4][250]  ( .E(n3586), .D(\vrf/N270 ), .Q(
        \vrf/regTable[4][250] ) );
  LHQD1BWP \vrf/regTable_reg[4][251]  ( .E(\vrf/N284 ), .D(\vrf/N271 ), .Q(
        \vrf/regTable[4][251] ) );
  LHQD1BWP \vrf/regTable_reg[4][252]  ( .E(n3586), .D(\vrf/N272 ), .Q(
        \vrf/regTable[4][252] ) );
  LHQD1BWP \vrf/regTable_reg[4][253]  ( .E(n3586), .D(\vrf/N273 ), .Q(
        \vrf/regTable[4][253] ) );
  LHQD1BWP \vrf/regTable_reg[4][254]  ( .E(n3586), .D(\vrf/N274 ), .Q(
        \vrf/regTable[4][254] ) );
  LHQD1BWP \vrf/regTable_reg[4][255]  ( .E(n3586), .D(\vrf/N275 ), .Q(
        \vrf/regTable[4][255] ) );
  LHQD1BWP \vrf/regTable_reg[3][0]  ( .E(n3587), .D(\vrf/N18 ), .Q(
        \vrf/regTable[3][0] ) );
  LHQD1BWP \vrf/regTable_reg[3][1]  ( .E(n3587), .D(\vrf/N19 ), .Q(
        \vrf/regTable[3][1] ) );
  LHQD1BWP \vrf/regTable_reg[3][2]  ( .E(n3587), .D(\vrf/N20 ), .Q(
        \vrf/regTable[3][2] ) );
  LHQD1BWP \vrf/regTable_reg[3][3]  ( .E(n3587), .D(\vrf/N21 ), .Q(
        \vrf/regTable[3][3] ) );
  LHQD1BWP \vrf/regTable_reg[3][4]  ( .E(n3587), .D(\vrf/N22 ), .Q(
        \vrf/regTable[3][4] ) );
  LHQD1BWP \vrf/regTable_reg[3][5]  ( .E(n3587), .D(\vrf/N23 ), .Q(
        \vrf/regTable[3][5] ) );
  LHQD1BWP \vrf/regTable_reg[3][6]  ( .E(n3587), .D(\vrf/N24 ), .Q(
        \vrf/regTable[3][6] ) );
  LHQD1BWP \vrf/regTable_reg[3][7]  ( .E(n3587), .D(\vrf/N25 ), .Q(
        \vrf/regTable[3][7] ) );
  LHQD1BWP \vrf/regTable_reg[3][8]  ( .E(n3587), .D(\vrf/N26 ), .Q(
        \vrf/regTable[3][8] ) );
  LHQD1BWP \vrf/regTable_reg[3][9]  ( .E(n3587), .D(\vrf/N27 ), .Q(
        \vrf/regTable[3][9] ) );
  LHQD1BWP \vrf/regTable_reg[3][10]  ( .E(n3587), .D(\vrf/N28 ), .Q(
        \vrf/regTable[3][10] ) );
  LHQD1BWP \vrf/regTable_reg[3][11]  ( .E(n3587), .D(\vrf/N29 ), .Q(
        \vrf/regTable[3][11] ) );
  LHQD1BWP \vrf/regTable_reg[3][12]  ( .E(n3587), .D(\vrf/N30 ), .Q(
        \vrf/regTable[3][12] ) );
  LHQD1BWP \vrf/regTable_reg[3][13]  ( .E(n3587), .D(\vrf/N31 ), .Q(
        \vrf/regTable[3][13] ) );
  LHQD1BWP \vrf/regTable_reg[3][14]  ( .E(n3587), .D(\vrf/N32 ), .Q(
        \vrf/regTable[3][14] ) );
  LHQD1BWP \vrf/regTable_reg[3][15]  ( .E(n3587), .D(\vrf/N33 ), .Q(
        \vrf/regTable[3][15] ) );
  LHQD1BWP \vrf/regTable_reg[3][16]  ( .E(n3587), .D(\vrf/N34 ), .Q(
        \vrf/regTable[3][16] ) );
  LHQD1BWP \vrf/regTable_reg[3][17]  ( .E(n3587), .D(\vrf/N35 ), .Q(
        \vrf/regTable[3][17] ) );
  LHQD1BWP \vrf/regTable_reg[3][18]  ( .E(n3587), .D(\vrf/N36 ), .Q(
        \vrf/regTable[3][18] ) );
  LHQD1BWP \vrf/regTable_reg[3][19]  ( .E(n3587), .D(\vrf/N37 ), .Q(
        \vrf/regTable[3][19] ) );
  LHQD1BWP \vrf/regTable_reg[3][20]  ( .E(n3587), .D(\vrf/N38 ), .Q(
        \vrf/regTable[3][20] ) );
  LHQD1BWP \vrf/regTable_reg[3][21]  ( .E(n3587), .D(\vrf/N39 ), .Q(
        \vrf/regTable[3][21] ) );
  LHQD1BWP \vrf/regTable_reg[3][22]  ( .E(n3587), .D(\vrf/N40 ), .Q(
        \vrf/regTable[3][22] ) );
  LHQD1BWP \vrf/regTable_reg[3][23]  ( .E(n3587), .D(\vrf/N41 ), .Q(
        \vrf/regTable[3][23] ) );
  LHQD1BWP \vrf/regTable_reg[3][24]  ( .E(n3587), .D(\vrf/N42 ), .Q(
        \vrf/regTable[3][24] ) );
  LHQD1BWP \vrf/regTable_reg[3][25]  ( .E(n3587), .D(\vrf/N43 ), .Q(
        \vrf/regTable[3][25] ) );
  LHQD1BWP \vrf/regTable_reg[3][26]  ( .E(n3587), .D(\vrf/N44 ), .Q(
        \vrf/regTable[3][26] ) );
  LHQD1BWP \vrf/regTable_reg[3][27]  ( .E(n3587), .D(\vrf/N45 ), .Q(
        \vrf/regTable[3][27] ) );
  LHQD1BWP \vrf/regTable_reg[3][28]  ( .E(n3587), .D(\vrf/N46 ), .Q(
        \vrf/regTable[3][28] ) );
  LHQD1BWP \vrf/regTable_reg[3][29]  ( .E(n3587), .D(\vrf/N47 ), .Q(
        \vrf/regTable[3][29] ) );
  LHQD1BWP \vrf/regTable_reg[3][30]  ( .E(n3587), .D(\vrf/N48 ), .Q(
        \vrf/regTable[3][30] ) );
  LHQD1BWP \vrf/regTable_reg[3][31]  ( .E(n3587), .D(\vrf/N49 ), .Q(
        \vrf/regTable[3][31] ) );
  LHQD1BWP \vrf/regTable_reg[3][32]  ( .E(n3587), .D(\vrf/N50 ), .Q(
        \vrf/regTable[3][32] ) );
  LHQD1BWP \vrf/regTable_reg[3][33]  ( .E(n3587), .D(\vrf/N51 ), .Q(
        \vrf/regTable[3][33] ) );
  LHQD1BWP \vrf/regTable_reg[3][34]  ( .E(n3587), .D(\vrf/N52 ), .Q(
        \vrf/regTable[3][34] ) );
  LHQD1BWP \vrf/regTable_reg[3][35]  ( .E(n3587), .D(\vrf/N53 ), .Q(
        \vrf/regTable[3][35] ) );
  LHQD1BWP \vrf/regTable_reg[3][36]  ( .E(n3587), .D(\vrf/N54 ), .Q(
        \vrf/regTable[3][36] ) );
  LHQD1BWP \vrf/regTable_reg[3][37]  ( .E(n3587), .D(\vrf/N55 ), .Q(
        \vrf/regTable[3][37] ) );
  LHQD1BWP \vrf/regTable_reg[3][38]  ( .E(n3587), .D(\vrf/N56 ), .Q(
        \vrf/regTable[3][38] ) );
  LHQD1BWP \vrf/regTable_reg[3][39]  ( .E(n3587), .D(\vrf/N57 ), .Q(
        \vrf/regTable[3][39] ) );
  LHQD1BWP \vrf/regTable_reg[3][40]  ( .E(n3587), .D(\vrf/N58 ), .Q(
        \vrf/regTable[3][40] ) );
  LHQD1BWP \vrf/regTable_reg[3][41]  ( .E(n3587), .D(\vrf/N59 ), .Q(
        \vrf/regTable[3][41] ) );
  LHQD1BWP \vrf/regTable_reg[3][42]  ( .E(n3587), .D(\vrf/N60 ), .Q(
        \vrf/regTable[3][42] ) );
  LHQD1BWP \vrf/regTable_reg[3][43]  ( .E(n3587), .D(\vrf/N61 ), .Q(
        \vrf/regTable[3][43] ) );
  LHQD1BWP \vrf/regTable_reg[3][44]  ( .E(n3587), .D(\vrf/N62 ), .Q(
        \vrf/regTable[3][44] ) );
  LHQD1BWP \vrf/regTable_reg[3][45]  ( .E(n3587), .D(\vrf/N63 ), .Q(
        \vrf/regTable[3][45] ) );
  LHQD1BWP \vrf/regTable_reg[3][46]  ( .E(n3587), .D(\vrf/N64 ), .Q(
        \vrf/regTable[3][46] ) );
  LHQD1BWP \vrf/regTable_reg[3][47]  ( .E(n3587), .D(\vrf/N65 ), .Q(
        \vrf/regTable[3][47] ) );
  LHQD1BWP \vrf/regTable_reg[3][48]  ( .E(n3587), .D(\vrf/N66 ), .Q(
        \vrf/regTable[3][48] ) );
  LHQD1BWP \vrf/regTable_reg[3][49]  ( .E(n3587), .D(\vrf/N67 ), .Q(
        \vrf/regTable[3][49] ) );
  LHQD1BWP \vrf/regTable_reg[3][50]  ( .E(n3587), .D(\vrf/N68 ), .Q(
        \vrf/regTable[3][50] ) );
  LHQD1BWP \vrf/regTable_reg[3][51]  ( .E(n3587), .D(\vrf/N69 ), .Q(
        \vrf/regTable[3][51] ) );
  LHQD1BWP \vrf/regTable_reg[3][52]  ( .E(n3587), .D(\vrf/N70 ), .Q(
        \vrf/regTable[3][52] ) );
  LHQD1BWP \vrf/regTable_reg[3][53]  ( .E(n3587), .D(\vrf/N71 ), .Q(
        \vrf/regTable[3][53] ) );
  LHQD1BWP \vrf/regTable_reg[3][54]  ( .E(n3587), .D(\vrf/N72 ), .Q(
        \vrf/regTable[3][54] ) );
  LHQD1BWP \vrf/regTable_reg[3][55]  ( .E(n3587), .D(\vrf/N73 ), .Q(
        \vrf/regTable[3][55] ) );
  LHQD1BWP \vrf/regTable_reg[3][56]  ( .E(n3587), .D(\vrf/N74 ), .Q(
        \vrf/regTable[3][56] ) );
  LHQD1BWP \vrf/regTable_reg[3][57]  ( .E(n3587), .D(\vrf/N75 ), .Q(
        \vrf/regTable[3][57] ) );
  LHQD1BWP \vrf/regTable_reg[3][58]  ( .E(n3587), .D(\vrf/N76 ), .Q(
        \vrf/regTable[3][58] ) );
  LHQD1BWP \vrf/regTable_reg[3][59]  ( .E(n3587), .D(\vrf/N77 ), .Q(
        \vrf/regTable[3][59] ) );
  LHQD1BWP \vrf/regTable_reg[3][60]  ( .E(n3587), .D(\vrf/N78 ), .Q(
        \vrf/regTable[3][60] ) );
  LHQD1BWP \vrf/regTable_reg[3][61]  ( .E(n3587), .D(\vrf/N79 ), .Q(
        \vrf/regTable[3][61] ) );
  LHQD1BWP \vrf/regTable_reg[3][62]  ( .E(n3587), .D(\vrf/N80 ), .Q(
        \vrf/regTable[3][62] ) );
  LHQD1BWP \vrf/regTable_reg[3][63]  ( .E(n3587), .D(\vrf/N81 ), .Q(
        \vrf/regTable[3][63] ) );
  LHQD1BWP \vrf/regTable_reg[3][64]  ( .E(n3587), .D(\vrf/N82 ), .Q(
        \vrf/regTable[3][64] ) );
  LHQD1BWP \vrf/regTable_reg[3][65]  ( .E(n3587), .D(\vrf/N83 ), .Q(
        \vrf/regTable[3][65] ) );
  LHQD1BWP \vrf/regTable_reg[3][66]  ( .E(n3587), .D(\vrf/N84 ), .Q(
        \vrf/regTable[3][66] ) );
  LHQD1BWP \vrf/regTable_reg[3][67]  ( .E(n3587), .D(\vrf/N85 ), .Q(
        \vrf/regTable[3][67] ) );
  LHQD1BWP \vrf/regTable_reg[3][68]  ( .E(n3587), .D(\vrf/N86 ), .Q(
        \vrf/regTable[3][68] ) );
  LHQD1BWP \vrf/regTable_reg[3][69]  ( .E(n3587), .D(\vrf/N87 ), .Q(
        \vrf/regTable[3][69] ) );
  LHQD1BWP \vrf/regTable_reg[3][70]  ( .E(n3587), .D(\vrf/N88 ), .Q(
        \vrf/regTable[3][70] ) );
  LHQD1BWP \vrf/regTable_reg[3][71]  ( .E(n3587), .D(\vrf/N89 ), .Q(
        \vrf/regTable[3][71] ) );
  LHQD1BWP \vrf/regTable_reg[3][72]  ( .E(n3587), .D(\vrf/N90 ), .Q(
        \vrf/regTable[3][72] ) );
  LHQD1BWP \vrf/regTable_reg[3][73]  ( .E(n3587), .D(\vrf/N91 ), .Q(
        \vrf/regTable[3][73] ) );
  LHQD1BWP \vrf/regTable_reg[3][74]  ( .E(n3587), .D(\vrf/N92 ), .Q(
        \vrf/regTable[3][74] ) );
  LHQD1BWP \vrf/regTable_reg[3][75]  ( .E(n3587), .D(\vrf/N93 ), .Q(
        \vrf/regTable[3][75] ) );
  LHQD1BWP \vrf/regTable_reg[3][76]  ( .E(n3587), .D(\vrf/N94 ), .Q(
        \vrf/regTable[3][76] ) );
  LHQD1BWP \vrf/regTable_reg[3][77]  ( .E(n3587), .D(\vrf/N95 ), .Q(
        \vrf/regTable[3][77] ) );
  LHQD1BWP \vrf/regTable_reg[3][78]  ( .E(n3587), .D(\vrf/N96 ), .Q(
        \vrf/regTable[3][78] ) );
  LHQD1BWP \vrf/regTable_reg[3][79]  ( .E(n3587), .D(\vrf/N97 ), .Q(
        \vrf/regTable[3][79] ) );
  LHQD1BWP \vrf/regTable_reg[3][80]  ( .E(n3587), .D(\vrf/N98 ), .Q(
        \vrf/regTable[3][80] ) );
  LHQD1BWP \vrf/regTable_reg[3][81]  ( .E(n3587), .D(\vrf/N99 ), .Q(
        \vrf/regTable[3][81] ) );
  LHQD1BWP \vrf/regTable_reg[3][82]  ( .E(n3587), .D(\vrf/N100 ), .Q(
        \vrf/regTable[3][82] ) );
  LHQD1BWP \vrf/regTable_reg[3][83]  ( .E(n3587), .D(\vrf/N101 ), .Q(
        \vrf/regTable[3][83] ) );
  LHQD1BWP \vrf/regTable_reg[3][84]  ( .E(n3587), .D(\vrf/N102 ), .Q(
        \vrf/regTable[3][84] ) );
  LHQD1BWP \vrf/regTable_reg[3][85]  ( .E(n3587), .D(\vrf/N103 ), .Q(
        \vrf/regTable[3][85] ) );
  LHQD1BWP \vrf/regTable_reg[3][86]  ( .E(n3587), .D(\vrf/N104 ), .Q(
        \vrf/regTable[3][86] ) );
  LHQD1BWP \vrf/regTable_reg[3][87]  ( .E(n3587), .D(\vrf/N105 ), .Q(
        \vrf/regTable[3][87] ) );
  LHQD1BWP \vrf/regTable_reg[3][88]  ( .E(n3587), .D(\vrf/N106 ), .Q(
        \vrf/regTable[3][88] ) );
  LHQD1BWP \vrf/regTable_reg[3][89]  ( .E(n3587), .D(\vrf/N107 ), .Q(
        \vrf/regTable[3][89] ) );
  LHQD1BWP \vrf/regTable_reg[3][90]  ( .E(n3587), .D(\vrf/N108 ), .Q(
        \vrf/regTable[3][90] ) );
  LHQD1BWP \vrf/regTable_reg[3][91]  ( .E(n3587), .D(\vrf/N109 ), .Q(
        \vrf/regTable[3][91] ) );
  LHQD1BWP \vrf/regTable_reg[3][92]  ( .E(n3587), .D(\vrf/N110 ), .Q(
        \vrf/regTable[3][92] ) );
  LHQD1BWP \vrf/regTable_reg[3][93]  ( .E(n3587), .D(\vrf/N111 ), .Q(
        \vrf/regTable[3][93] ) );
  LHQD1BWP \vrf/regTable_reg[3][94]  ( .E(n3587), .D(\vrf/N112 ), .Q(
        \vrf/regTable[3][94] ) );
  LHQD1BWP \vrf/regTable_reg[3][95]  ( .E(n3587), .D(\vrf/N113 ), .Q(
        \vrf/regTable[3][95] ) );
  LHQD1BWP \vrf/regTable_reg[3][96]  ( .E(n3587), .D(\vrf/N114 ), .Q(
        \vrf/regTable[3][96] ) );
  LHQD1BWP \vrf/regTable_reg[3][97]  ( .E(n3587), .D(\vrf/N115 ), .Q(
        \vrf/regTable[3][97] ) );
  LHQD1BWP \vrf/regTable_reg[3][98]  ( .E(n3587), .D(\vrf/N116 ), .Q(
        \vrf/regTable[3][98] ) );
  LHQD1BWP \vrf/regTable_reg[3][99]  ( .E(n3587), .D(\vrf/N118 ), .Q(
        \vrf/regTable[3][99] ) );
  LHQD1BWP \vrf/regTable_reg[3][100]  ( .E(n3587), .D(\vrf/N119 ), .Q(
        \vrf/regTable[3][100] ) );
  LHQD1BWP \vrf/regTable_reg[3][101]  ( .E(n3587), .D(\vrf/N120 ), .Q(
        \vrf/regTable[3][101] ) );
  LHQD1BWP \vrf/regTable_reg[3][102]  ( .E(n3587), .D(\vrf/N121 ), .Q(
        \vrf/regTable[3][102] ) );
  LHQD1BWP \vrf/regTable_reg[3][103]  ( .E(n3587), .D(\vrf/N122 ), .Q(
        \vrf/regTable[3][103] ) );
  LHQD1BWP \vrf/regTable_reg[3][104]  ( .E(n3587), .D(\vrf/N123 ), .Q(
        \vrf/regTable[3][104] ) );
  LHQD1BWP \vrf/regTable_reg[3][105]  ( .E(n3587), .D(\vrf/N124 ), .Q(
        \vrf/regTable[3][105] ) );
  LHQD1BWP \vrf/regTable_reg[3][106]  ( .E(n3587), .D(\vrf/N125 ), .Q(
        \vrf/regTable[3][106] ) );
  LHQD1BWP \vrf/regTable_reg[3][107]  ( .E(n3587), .D(\vrf/N126 ), .Q(
        \vrf/regTable[3][107] ) );
  LHQD1BWP \vrf/regTable_reg[3][108]  ( .E(n3587), .D(\vrf/N127 ), .Q(
        \vrf/regTable[3][108] ) );
  LHQD1BWP \vrf/regTable_reg[3][109]  ( .E(n3587), .D(\vrf/N128 ), .Q(
        \vrf/regTable[3][109] ) );
  LHQD1BWP \vrf/regTable_reg[3][110]  ( .E(n3587), .D(\vrf/N129 ), .Q(
        \vrf/regTable[3][110] ) );
  LHQD1BWP \vrf/regTable_reg[3][111]  ( .E(n3587), .D(\vrf/N130 ), .Q(
        \vrf/regTable[3][111] ) );
  LHQD1BWP \vrf/regTable_reg[3][112]  ( .E(n3587), .D(\vrf/N131 ), .Q(
        \vrf/regTable[3][112] ) );
  LHQD1BWP \vrf/regTable_reg[3][113]  ( .E(n3587), .D(\vrf/N132 ), .Q(
        \vrf/regTable[3][113] ) );
  LHQD1BWP \vrf/regTable_reg[3][114]  ( .E(n3587), .D(\vrf/N133 ), .Q(
        \vrf/regTable[3][114] ) );
  LHQD1BWP \vrf/regTable_reg[3][115]  ( .E(n3587), .D(\vrf/N134 ), .Q(
        \vrf/regTable[3][115] ) );
  LHQD1BWP \vrf/regTable_reg[3][116]  ( .E(n3587), .D(\vrf/N135 ), .Q(
        \vrf/regTable[3][116] ) );
  LHQD1BWP \vrf/regTable_reg[3][117]  ( .E(n3587), .D(\vrf/N136 ), .Q(
        \vrf/regTable[3][117] ) );
  LHQD1BWP \vrf/regTable_reg[3][118]  ( .E(n3587), .D(\vrf/N137 ), .Q(
        \vrf/regTable[3][118] ) );
  LHQD1BWP \vrf/regTable_reg[3][119]  ( .E(n3587), .D(\vrf/N138 ), .Q(
        \vrf/regTable[3][119] ) );
  LHQD1BWP \vrf/regTable_reg[3][120]  ( .E(n3587), .D(\vrf/N139 ), .Q(
        \vrf/regTable[3][120] ) );
  LHQD1BWP \vrf/regTable_reg[3][121]  ( .E(n3587), .D(\vrf/N140 ), .Q(
        \vrf/regTable[3][121] ) );
  LHQD1BWP \vrf/regTable_reg[3][122]  ( .E(n3587), .D(\vrf/N141 ), .Q(
        \vrf/regTable[3][122] ) );
  LHQD1BWP \vrf/regTable_reg[3][123]  ( .E(n3587), .D(\vrf/N142 ), .Q(
        \vrf/regTable[3][123] ) );
  LHQD1BWP \vrf/regTable_reg[3][124]  ( .E(n3587), .D(\vrf/N143 ), .Q(
        \vrf/regTable[3][124] ) );
  LHQD1BWP \vrf/regTable_reg[3][125]  ( .E(n3587), .D(\vrf/N144 ), .Q(
        \vrf/regTable[3][125] ) );
  LHQD1BWP \vrf/regTable_reg[3][126]  ( .E(n3587), .D(\vrf/N145 ), .Q(
        \vrf/regTable[3][126] ) );
  LHQD1BWP \vrf/regTable_reg[3][127]  ( .E(n3587), .D(\vrf/N146 ), .Q(
        \vrf/regTable[3][127] ) );
  LHQD1BWP \vrf/regTable_reg[3][128]  ( .E(n3587), .D(\vrf/N147 ), .Q(
        \vrf/regTable[3][128] ) );
  LHQD1BWP \vrf/regTable_reg[3][129]  ( .E(n3587), .D(\vrf/N148 ), .Q(
        \vrf/regTable[3][129] ) );
  LHQD1BWP \vrf/regTable_reg[3][130]  ( .E(n3587), .D(\vrf/N149 ), .Q(
        \vrf/regTable[3][130] ) );
  LHQD1BWP \vrf/regTable_reg[3][131]  ( .E(n3587), .D(\vrf/N150 ), .Q(
        \vrf/regTable[3][131] ) );
  LHQD1BWP \vrf/regTable_reg[3][132]  ( .E(n3587), .D(\vrf/N151 ), .Q(
        \vrf/regTable[3][132] ) );
  LHQD1BWP \vrf/regTable_reg[3][133]  ( .E(n3587), .D(\vrf/N152 ), .Q(
        \vrf/regTable[3][133] ) );
  LHQD1BWP \vrf/regTable_reg[3][134]  ( .E(n3587), .D(\vrf/N153 ), .Q(
        \vrf/regTable[3][134] ) );
  LHQD1BWP \vrf/regTable_reg[3][135]  ( .E(n3587), .D(\vrf/N154 ), .Q(
        \vrf/regTable[3][135] ) );
  LHQD1BWP \vrf/regTable_reg[3][136]  ( .E(n3587), .D(\vrf/N155 ), .Q(
        \vrf/regTable[3][136] ) );
  LHQD1BWP \vrf/regTable_reg[3][137]  ( .E(\vrf/N287 ), .D(\vrf/N156 ), .Q(
        \vrf/regTable[3][137] ) );
  LHQD1BWP \vrf/regTable_reg[3][138]  ( .E(n3587), .D(\vrf/N157 ), .Q(
        \vrf/regTable[3][138] ) );
  LHQD1BWP \vrf/regTable_reg[3][139]  ( .E(\vrf/N287 ), .D(\vrf/N158 ), .Q(
        \vrf/regTable[3][139] ) );
  LHQD1BWP \vrf/regTable_reg[3][140]  ( .E(n3587), .D(\vrf/N159 ), .Q(
        \vrf/regTable[3][140] ) );
  LHQD1BWP \vrf/regTable_reg[3][141]  ( .E(\vrf/N287 ), .D(\vrf/N160 ), .Q(
        \vrf/regTable[3][141] ) );
  LHQD1BWP \vrf/regTable_reg[3][142]  ( .E(n3587), .D(\vrf/N161 ), .Q(
        \vrf/regTable[3][142] ) );
  LHQD1BWP \vrf/regTable_reg[3][143]  ( .E(\vrf/N287 ), .D(\vrf/N162 ), .Q(
        \vrf/regTable[3][143] ) );
  LHQD1BWP \vrf/regTable_reg[3][144]  ( .E(n3587), .D(\vrf/N163 ), .Q(
        \vrf/regTable[3][144] ) );
  LHQD1BWP \vrf/regTable_reg[3][145]  ( .E(\vrf/N287 ), .D(\vrf/N164 ), .Q(
        \vrf/regTable[3][145] ) );
  LHQD1BWP \vrf/regTable_reg[3][146]  ( .E(n3587), .D(\vrf/N165 ), .Q(
        \vrf/regTable[3][146] ) );
  LHQD1BWP \vrf/regTable_reg[3][147]  ( .E(\vrf/N287 ), .D(\vrf/N166 ), .Q(
        \vrf/regTable[3][147] ) );
  LHQD1BWP \vrf/regTable_reg[3][148]  ( .E(n3587), .D(\vrf/N167 ), .Q(
        \vrf/regTable[3][148] ) );
  LHQD1BWP \vrf/regTable_reg[3][149]  ( .E(n3587), .D(\vrf/N168 ), .Q(
        \vrf/regTable[3][149] ) );
  LHQD1BWP \vrf/regTable_reg[3][150]  ( .E(n3587), .D(\vrf/N169 ), .Q(
        \vrf/regTable[3][150] ) );
  LHQD1BWP \vrf/regTable_reg[3][151]  ( .E(\vrf/N287 ), .D(\vrf/N170 ), .Q(
        \vrf/regTable[3][151] ) );
  LHQD1BWP \vrf/regTable_reg[3][152]  ( .E(n3587), .D(\vrf/N171 ), .Q(
        \vrf/regTable[3][152] ) );
  LHQD1BWP \vrf/regTable_reg[3][153]  ( .E(n3587), .D(\vrf/N172 ), .Q(
        \vrf/regTable[3][153] ) );
  LHQD1BWP \vrf/regTable_reg[3][154]  ( .E(n3587), .D(\vrf/N173 ), .Q(
        \vrf/regTable[3][154] ) );
  LHQD1BWP \vrf/regTable_reg[3][155]  ( .E(\vrf/N287 ), .D(\vrf/N174 ), .Q(
        \vrf/regTable[3][155] ) );
  LHQD1BWP \vrf/regTable_reg[3][156]  ( .E(n3587), .D(\vrf/N175 ), .Q(
        \vrf/regTable[3][156] ) );
  LHQD1BWP \vrf/regTable_reg[3][157]  ( .E(n3587), .D(\vrf/N176 ), .Q(
        \vrf/regTable[3][157] ) );
  LHQD1BWP \vrf/regTable_reg[3][158]  ( .E(n3587), .D(\vrf/N177 ), .Q(
        \vrf/regTable[3][158] ) );
  LHQD1BWP \vrf/regTable_reg[3][159]  ( .E(n3587), .D(\vrf/N178 ), .Q(
        \vrf/regTable[3][159] ) );
  LHQD1BWP \vrf/regTable_reg[3][160]  ( .E(\vrf/N287 ), .D(\vrf/N179 ), .Q(
        \vrf/regTable[3][160] ) );
  LHQD1BWP \vrf/regTable_reg[3][161]  ( .E(n3587), .D(\vrf/N180 ), .Q(
        \vrf/regTable[3][161] ) );
  LHQD1BWP \vrf/regTable_reg[3][162]  ( .E(n3587), .D(\vrf/N181 ), .Q(
        \vrf/regTable[3][162] ) );
  LHQD1BWP \vrf/regTable_reg[3][163]  ( .E(n3587), .D(\vrf/N182 ), .Q(
        \vrf/regTable[3][163] ) );
  LHQD1BWP \vrf/regTable_reg[3][164]  ( .E(\vrf/N287 ), .D(\vrf/N183 ), .Q(
        \vrf/regTable[3][164] ) );
  LHQD1BWP \vrf/regTable_reg[3][165]  ( .E(n3587), .D(\vrf/N184 ), .Q(
        \vrf/regTable[3][165] ) );
  LHQD1BWP \vrf/regTable_reg[3][166]  ( .E(n3587), .D(\vrf/N185 ), .Q(
        \vrf/regTable[3][166] ) );
  LHQD1BWP \vrf/regTable_reg[3][167]  ( .E(n3587), .D(\vrf/N186 ), .Q(
        \vrf/regTable[3][167] ) );
  LHQD1BWP \vrf/regTable_reg[3][168]  ( .E(\vrf/N287 ), .D(\vrf/N187 ), .Q(
        \vrf/regTable[3][168] ) );
  LHQD1BWP \vrf/regTable_reg[3][169]  ( .E(n3587), .D(\vrf/N188 ), .Q(
        \vrf/regTable[3][169] ) );
  LHQD1BWP \vrf/regTable_reg[3][170]  ( .E(n3587), .D(\vrf/N189 ), .Q(
        \vrf/regTable[3][170] ) );
  LHQD1BWP \vrf/regTable_reg[3][171]  ( .E(n3587), .D(\vrf/N190 ), .Q(
        \vrf/regTable[3][171] ) );
  LHQD1BWP \vrf/regTable_reg[3][172]  ( .E(n3587), .D(\vrf/N191 ), .Q(
        \vrf/regTable[3][172] ) );
  LHQD1BWP \vrf/regTable_reg[3][173]  ( .E(n3587), .D(\vrf/N192 ), .Q(
        \vrf/regTable[3][173] ) );
  LHQD1BWP \vrf/regTable_reg[3][174]  ( .E(\vrf/N287 ), .D(\vrf/N193 ), .Q(
        \vrf/regTable[3][174] ) );
  LHQD1BWP \vrf/regTable_reg[3][175]  ( .E(n3587), .D(\vrf/N194 ), .Q(
        \vrf/regTable[3][175] ) );
  LHQD1BWP \vrf/regTable_reg[3][176]  ( .E(n3587), .D(\vrf/N195 ), .Q(
        \vrf/regTable[3][176] ) );
  LHQD1BWP \vrf/regTable_reg[3][177]  ( .E(n3587), .D(\vrf/N196 ), .Q(
        \vrf/regTable[3][177] ) );
  LHQD1BWP \vrf/regTable_reg[3][178]  ( .E(n3587), .D(\vrf/N197 ), .Q(
        \vrf/regTable[3][178] ) );
  LHQD1BWP \vrf/regTable_reg[3][179]  ( .E(\vrf/N287 ), .D(\vrf/N198 ), .Q(
        \vrf/regTable[3][179] ) );
  LHQD1BWP \vrf/regTable_reg[3][180]  ( .E(n3587), .D(\vrf/N199 ), .Q(
        \vrf/regTable[3][180] ) );
  LHQD1BWP \vrf/regTable_reg[3][181]  ( .E(n3587), .D(\vrf/N200 ), .Q(
        \vrf/regTable[3][181] ) );
  LHQD1BWP \vrf/regTable_reg[3][182]  ( .E(n3587), .D(\vrf/N201 ), .Q(
        \vrf/regTable[3][182] ) );
  LHQD1BWP \vrf/regTable_reg[3][183]  ( .E(n3587), .D(\vrf/N202 ), .Q(
        \vrf/regTable[3][183] ) );
  LHQD1BWP \vrf/regTable_reg[3][184]  ( .E(n3587), .D(\vrf/N203 ), .Q(
        \vrf/regTable[3][184] ) );
  LHQD1BWP \vrf/regTable_reg[3][185]  ( .E(n3587), .D(\vrf/N204 ), .Q(
        \vrf/regTable[3][185] ) );
  LHQD1BWP \vrf/regTable_reg[3][186]  ( .E(n3587), .D(\vrf/N205 ), .Q(
        \vrf/regTable[3][186] ) );
  LHQD1BWP \vrf/regTable_reg[3][187]  ( .E(n3587), .D(\vrf/N206 ), .Q(
        \vrf/regTable[3][187] ) );
  LHQD1BWP \vrf/regTable_reg[3][188]  ( .E(n3587), .D(\vrf/N207 ), .Q(
        \vrf/regTable[3][188] ) );
  LHQD1BWP \vrf/regTable_reg[3][189]  ( .E(\vrf/N287 ), .D(\vrf/N208 ), .Q(
        \vrf/regTable[3][189] ) );
  LHQD1BWP \vrf/regTable_reg[3][190]  ( .E(n3587), .D(\vrf/N209 ), .Q(
        \vrf/regTable[3][190] ) );
  LHQD1BWP \vrf/regTable_reg[3][191]  ( .E(n3587), .D(\vrf/N210 ), .Q(
        \vrf/regTable[3][191] ) );
  LHQD1BWP \vrf/regTable_reg[3][192]  ( .E(n3587), .D(\vrf/N211 ), .Q(
        \vrf/regTable[3][192] ) );
  LHQD1BWP \vrf/regTable_reg[3][193]  ( .E(n3587), .D(\vrf/N212 ), .Q(
        \vrf/regTable[3][193] ) );
  LHQD1BWP \vrf/regTable_reg[3][194]  ( .E(\vrf/N287 ), .D(\vrf/N213 ), .Q(
        \vrf/regTable[3][194] ) );
  LHQD1BWP \vrf/regTable_reg[3][195]  ( .E(\vrf/N287 ), .D(\vrf/N214 ), .Q(
        \vrf/regTable[3][195] ) );
  LHQD1BWP \vrf/regTable_reg[3][196]  ( .E(n3587), .D(\vrf/N215 ), .Q(
        \vrf/regTable[3][196] ) );
  LHQD1BWP \vrf/regTable_reg[3][197]  ( .E(n3587), .D(\vrf/N216 ), .Q(
        \vrf/regTable[3][197] ) );
  LHQD1BWP \vrf/regTable_reg[3][198]  ( .E(n3587), .D(\vrf/N218 ), .Q(
        \vrf/regTable[3][198] ) );
  LHQD1BWP \vrf/regTable_reg[3][199]  ( .E(n3587), .D(\vrf/N219 ), .Q(
        \vrf/regTable[3][199] ) );
  LHQD1BWP \vrf/regTable_reg[3][200]  ( .E(n3587), .D(\vrf/N220 ), .Q(
        \vrf/regTable[3][200] ) );
  LHQD1BWP \vrf/regTable_reg[3][201]  ( .E(\vrf/N287 ), .D(\vrf/N221 ), .Q(
        \vrf/regTable[3][201] ) );
  LHQD1BWP \vrf/regTable_reg[3][202]  ( .E(n3587), .D(\vrf/N222 ), .Q(
        \vrf/regTable[3][202] ) );
  LHQD1BWP \vrf/regTable_reg[3][203]  ( .E(n3587), .D(\vrf/N223 ), .Q(
        \vrf/regTable[3][203] ) );
  LHQD1BWP \vrf/regTable_reg[3][204]  ( .E(\vrf/N287 ), .D(\vrf/N224 ), .Q(
        \vrf/regTable[3][204] ) );
  LHQD1BWP \vrf/regTable_reg[3][205]  ( .E(n3587), .D(\vrf/N225 ), .Q(
        \vrf/regTable[3][205] ) );
  LHQD1BWP \vrf/regTable_reg[3][206]  ( .E(\vrf/N287 ), .D(\vrf/N226 ), .Q(
        \vrf/regTable[3][206] ) );
  LHQD1BWP \vrf/regTable_reg[3][207]  ( .E(n3587), .D(\vrf/N227 ), .Q(
        \vrf/regTable[3][207] ) );
  LHQD1BWP \vrf/regTable_reg[3][208]  ( .E(n3587), .D(\vrf/N228 ), .Q(
        \vrf/regTable[3][208] ) );
  LHQD1BWP \vrf/regTable_reg[3][209]  ( .E(n3587), .D(\vrf/N229 ), .Q(
        \vrf/regTable[3][209] ) );
  LHQD1BWP \vrf/regTable_reg[3][210]  ( .E(n3587), .D(\vrf/N230 ), .Q(
        \vrf/regTable[3][210] ) );
  LHQD1BWP \vrf/regTable_reg[3][211]  ( .E(n3587), .D(\vrf/N231 ), .Q(
        \vrf/regTable[3][211] ) );
  LHQD1BWP \vrf/regTable_reg[3][212]  ( .E(n3587), .D(\vrf/N232 ), .Q(
        \vrf/regTable[3][212] ) );
  LHQD1BWP \vrf/regTable_reg[3][213]  ( .E(n3587), .D(\vrf/N233 ), .Q(
        \vrf/regTable[3][213] ) );
  LHQD1BWP \vrf/regTable_reg[3][214]  ( .E(n3587), .D(\vrf/N234 ), .Q(
        \vrf/regTable[3][214] ) );
  LHQD1BWP \vrf/regTable_reg[3][215]  ( .E(n3587), .D(\vrf/N235 ), .Q(
        \vrf/regTable[3][215] ) );
  LHQD1BWP \vrf/regTable_reg[3][216]  ( .E(n3587), .D(\vrf/N236 ), .Q(
        \vrf/regTable[3][216] ) );
  LHQD1BWP \vrf/regTable_reg[3][217]  ( .E(n3587), .D(\vrf/N237 ), .Q(
        \vrf/regTable[3][217] ) );
  LHQD1BWP \vrf/regTable_reg[3][218]  ( .E(n3587), .D(\vrf/N238 ), .Q(
        \vrf/regTable[3][218] ) );
  LHQD1BWP \vrf/regTable_reg[3][219]  ( .E(n3587), .D(\vrf/N239 ), .Q(
        \vrf/regTable[3][219] ) );
  LHQD1BWP \vrf/regTable_reg[3][220]  ( .E(n3587), .D(\vrf/N240 ), .Q(
        \vrf/regTable[3][220] ) );
  LHQD1BWP \vrf/regTable_reg[3][221]  ( .E(n3587), .D(\vrf/N241 ), .Q(
        \vrf/regTable[3][221] ) );
  LHQD1BWP \vrf/regTable_reg[3][222]  ( .E(n3587), .D(\vrf/N242 ), .Q(
        \vrf/regTable[3][222] ) );
  LHQD1BWP \vrf/regTable_reg[3][223]  ( .E(\vrf/N287 ), .D(\vrf/N243 ), .Q(
        \vrf/regTable[3][223] ) );
  LHQD1BWP \vrf/regTable_reg[3][224]  ( .E(n3587), .D(\vrf/N244 ), .Q(
        \vrf/regTable[3][224] ) );
  LHQD1BWP \vrf/regTable_reg[3][225]  ( .E(n3587), .D(\vrf/N245 ), .Q(
        \vrf/regTable[3][225] ) );
  LHQD1BWP \vrf/regTable_reg[3][226]  ( .E(n3587), .D(\vrf/N246 ), .Q(
        \vrf/regTable[3][226] ) );
  LHQD1BWP \vrf/regTable_reg[3][227]  ( .E(\vrf/N287 ), .D(\vrf/N247 ), .Q(
        \vrf/regTable[3][227] ) );
  LHQD1BWP \vrf/regTable_reg[3][228]  ( .E(n3587), .D(\vrf/N248 ), .Q(
        \vrf/regTable[3][228] ) );
  LHQD1BWP \vrf/regTable_reg[3][229]  ( .E(n3587), .D(\vrf/N249 ), .Q(
        \vrf/regTable[3][229] ) );
  LHQD1BWP \vrf/regTable_reg[3][230]  ( .E(n3587), .D(\vrf/N250 ), .Q(
        \vrf/regTable[3][230] ) );
  LHQD1BWP \vrf/regTable_reg[3][231]  ( .E(\vrf/N287 ), .D(\vrf/N251 ), .Q(
        \vrf/regTable[3][231] ) );
  LHQD1BWP \vrf/regTable_reg[3][232]  ( .E(n3587), .D(\vrf/N252 ), .Q(
        \vrf/regTable[3][232] ) );
  LHQD1BWP \vrf/regTable_reg[3][233]  ( .E(n3587), .D(\vrf/N253 ), .Q(
        \vrf/regTable[3][233] ) );
  LHQD1BWP \vrf/regTable_reg[3][234]  ( .E(n3587), .D(\vrf/N254 ), .Q(
        \vrf/regTable[3][234] ) );
  LHQD1BWP \vrf/regTable_reg[3][235]  ( .E(n3587), .D(\vrf/N255 ), .Q(
        \vrf/regTable[3][235] ) );
  LHQD1BWP \vrf/regTable_reg[3][236]  ( .E(n3587), .D(\vrf/N256 ), .Q(
        \vrf/regTable[3][236] ) );
  LHQD1BWP \vrf/regTable_reg[3][237]  ( .E(n3587), .D(\vrf/N257 ), .Q(
        \vrf/regTable[3][237] ) );
  LHQD1BWP \vrf/regTable_reg[3][238]  ( .E(n3587), .D(\vrf/N258 ), .Q(
        \vrf/regTable[3][238] ) );
  LHQD1BWP \vrf/regTable_reg[3][239]  ( .E(n3587), .D(\vrf/N259 ), .Q(
        \vrf/regTable[3][239] ) );
  LHQD1BWP \vrf/regTable_reg[3][240]  ( .E(n3587), .D(\vrf/N260 ), .Q(
        \vrf/regTable[3][240] ) );
  LHQD1BWP \vrf/regTable_reg[3][241]  ( .E(n3587), .D(\vrf/N261 ), .Q(
        \vrf/regTable[3][241] ) );
  LHQD1BWP \vrf/regTable_reg[3][242]  ( .E(n3587), .D(\vrf/N262 ), .Q(
        \vrf/regTable[3][242] ) );
  LHQD1BWP \vrf/regTable_reg[3][243]  ( .E(n3587), .D(\vrf/N263 ), .Q(
        \vrf/regTable[3][243] ) );
  LHQD1BWP \vrf/regTable_reg[3][244]  ( .E(n3587), .D(\vrf/N264 ), .Q(
        \vrf/regTable[3][244] ) );
  LHQD1BWP \vrf/regTable_reg[3][245]  ( .E(n3587), .D(\vrf/N265 ), .Q(
        \vrf/regTable[3][245] ) );
  LHQD1BWP \vrf/regTable_reg[3][246]  ( .E(n3587), .D(\vrf/N266 ), .Q(
        \vrf/regTable[3][246] ) );
  LHQD1BWP \vrf/regTable_reg[3][247]  ( .E(n3587), .D(\vrf/N267 ), .Q(
        \vrf/regTable[3][247] ) );
  LHQD1BWP \vrf/regTable_reg[3][248]  ( .E(n3587), .D(\vrf/N268 ), .Q(
        \vrf/regTable[3][248] ) );
  LHQD1BWP \vrf/regTable_reg[3][249]  ( .E(n3587), .D(\vrf/N269 ), .Q(
        \vrf/regTable[3][249] ) );
  LHQD1BWP \vrf/regTable_reg[3][250]  ( .E(n3587), .D(\vrf/N270 ), .Q(
        \vrf/regTable[3][250] ) );
  LHQD1BWP \vrf/regTable_reg[3][251]  ( .E(\vrf/N287 ), .D(\vrf/N271 ), .Q(
        \vrf/regTable[3][251] ) );
  LHQD1BWP \vrf/regTable_reg[3][252]  ( .E(n3587), .D(\vrf/N272 ), .Q(
        \vrf/regTable[3][252] ) );
  LHQD1BWP \vrf/regTable_reg[3][253]  ( .E(n3587), .D(\vrf/N273 ), .Q(
        \vrf/regTable[3][253] ) );
  LHQD1BWP \vrf/regTable_reg[3][254]  ( .E(n3587), .D(\vrf/N274 ), .Q(
        \vrf/regTable[3][254] ) );
  LHQD1BWP \vrf/regTable_reg[3][255]  ( .E(n3587), .D(\vrf/N275 ), .Q(
        \vrf/regTable[3][255] ) );
  LHQD1BWP \vrf/regTable_reg[2][0]  ( .E(n3589), .D(\vrf/N18 ), .Q(
        \vrf/regTable[2][0] ) );
  LHQD1BWP \vrf/regTable_reg[2][1]  ( .E(n3589), .D(\vrf/N19 ), .Q(
        \vrf/regTable[2][1] ) );
  LHQD1BWP \vrf/regTable_reg[2][2]  ( .E(n3589), .D(\vrf/N20 ), .Q(
        \vrf/regTable[2][2] ) );
  LHQD1BWP \vrf/regTable_reg[2][3]  ( .E(n3589), .D(\vrf/N21 ), .Q(
        \vrf/regTable[2][3] ) );
  LHQD1BWP \vrf/regTable_reg[2][4]  ( .E(n3589), .D(\vrf/N22 ), .Q(
        \vrf/regTable[2][4] ) );
  LHQD1BWP \vrf/regTable_reg[2][5]  ( .E(n3589), .D(\vrf/N23 ), .Q(
        \vrf/regTable[2][5] ) );
  LHQD1BWP \vrf/regTable_reg[2][6]  ( .E(n3589), .D(\vrf/N24 ), .Q(
        \vrf/regTable[2][6] ) );
  LHQD1BWP \vrf/regTable_reg[2][7]  ( .E(n3589), .D(\vrf/N25 ), .Q(
        \vrf/regTable[2][7] ) );
  LHQD1BWP \vrf/regTable_reg[2][8]  ( .E(n3589), .D(\vrf/N26 ), .Q(
        \vrf/regTable[2][8] ) );
  LHQD1BWP \vrf/regTable_reg[2][9]  ( .E(n3589), .D(\vrf/N27 ), .Q(
        \vrf/regTable[2][9] ) );
  LHQD1BWP \vrf/regTable_reg[2][10]  ( .E(n3589), .D(\vrf/N28 ), .Q(
        \vrf/regTable[2][10] ) );
  LHQD1BWP \vrf/regTable_reg[2][11]  ( .E(n3589), .D(\vrf/N29 ), .Q(
        \vrf/regTable[2][11] ) );
  LHQD1BWP \vrf/regTable_reg[2][12]  ( .E(n3589), .D(\vrf/N30 ), .Q(
        \vrf/regTable[2][12] ) );
  LHQD1BWP \vrf/regTable_reg[2][13]  ( .E(n3589), .D(\vrf/N31 ), .Q(
        \vrf/regTable[2][13] ) );
  LHQD1BWP \vrf/regTable_reg[2][14]  ( .E(n3589), .D(\vrf/N32 ), .Q(
        \vrf/regTable[2][14] ) );
  LHQD1BWP \vrf/regTable_reg[2][15]  ( .E(n3589), .D(\vrf/N33 ), .Q(
        \vrf/regTable[2][15] ) );
  LHQD1BWP \vrf/regTable_reg[2][16]  ( .E(n3589), .D(\vrf/N34 ), .Q(
        \vrf/regTable[2][16] ) );
  LHQD1BWP \vrf/regTable_reg[2][17]  ( .E(n3589), .D(\vrf/N35 ), .Q(
        \vrf/regTable[2][17] ) );
  LHQD1BWP \vrf/regTable_reg[2][18]  ( .E(n3589), .D(\vrf/N36 ), .Q(
        \vrf/regTable[2][18] ) );
  LHQD1BWP \vrf/regTable_reg[2][19]  ( .E(n3589), .D(\vrf/N37 ), .Q(
        \vrf/regTable[2][19] ) );
  LHQD1BWP \vrf/regTable_reg[2][20]  ( .E(n3589), .D(\vrf/N38 ), .Q(
        \vrf/regTable[2][20] ) );
  LHQD1BWP \vrf/regTable_reg[2][21]  ( .E(n3589), .D(\vrf/N39 ), .Q(
        \vrf/regTable[2][21] ) );
  LHQD1BWP \vrf/regTable_reg[2][22]  ( .E(n3589), .D(\vrf/N40 ), .Q(
        \vrf/regTable[2][22] ) );
  LHQD1BWP \vrf/regTable_reg[2][23]  ( .E(n3589), .D(\vrf/N41 ), .Q(
        \vrf/regTable[2][23] ) );
  LHQD1BWP \vrf/regTable_reg[2][24]  ( .E(n3589), .D(\vrf/N42 ), .Q(
        \vrf/regTable[2][24] ) );
  LHQD1BWP \vrf/regTable_reg[2][25]  ( .E(n3589), .D(\vrf/N43 ), .Q(
        \vrf/regTable[2][25] ) );
  LHQD1BWP \vrf/regTable_reg[2][26]  ( .E(n3589), .D(\vrf/N44 ), .Q(
        \vrf/regTable[2][26] ) );
  LHQD1BWP \vrf/regTable_reg[2][27]  ( .E(n3589), .D(\vrf/N45 ), .Q(
        \vrf/regTable[2][27] ) );
  LHQD1BWP \vrf/regTable_reg[2][28]  ( .E(n3589), .D(\vrf/N46 ), .Q(
        \vrf/regTable[2][28] ) );
  LHQD1BWP \vrf/regTable_reg[2][29]  ( .E(n3589), .D(\vrf/N47 ), .Q(
        \vrf/regTable[2][29] ) );
  LHQD1BWP \vrf/regTable_reg[2][30]  ( .E(n3589), .D(\vrf/N48 ), .Q(
        \vrf/regTable[2][30] ) );
  LHQD1BWP \vrf/regTable_reg[2][31]  ( .E(n3589), .D(\vrf/N49 ), .Q(
        \vrf/regTable[2][31] ) );
  LHQD1BWP \vrf/regTable_reg[2][32]  ( .E(n3589), .D(\vrf/N50 ), .Q(
        \vrf/regTable[2][32] ) );
  LHQD1BWP \vrf/regTable_reg[2][33]  ( .E(n3589), .D(\vrf/N51 ), .Q(
        \vrf/regTable[2][33] ) );
  LHQD1BWP \vrf/regTable_reg[2][34]  ( .E(n3589), .D(\vrf/N52 ), .Q(
        \vrf/regTable[2][34] ) );
  LHQD1BWP \vrf/regTable_reg[2][35]  ( .E(n3589), .D(\vrf/N53 ), .Q(
        \vrf/regTable[2][35] ) );
  LHQD1BWP \vrf/regTable_reg[2][36]  ( .E(n3589), .D(\vrf/N54 ), .Q(
        \vrf/regTable[2][36] ) );
  LHQD1BWP \vrf/regTable_reg[2][37]  ( .E(n3589), .D(\vrf/N55 ), .Q(
        \vrf/regTable[2][37] ) );
  LHQD1BWP \vrf/regTable_reg[2][38]  ( .E(n3589), .D(\vrf/N56 ), .Q(
        \vrf/regTable[2][38] ) );
  LHQD1BWP \vrf/regTable_reg[2][39]  ( .E(n3589), .D(\vrf/N57 ), .Q(
        \vrf/regTable[2][39] ) );
  LHQD1BWP \vrf/regTable_reg[2][40]  ( .E(n3589), .D(\vrf/N58 ), .Q(
        \vrf/regTable[2][40] ) );
  LHQD1BWP \vrf/regTable_reg[2][41]  ( .E(n3589), .D(\vrf/N59 ), .Q(
        \vrf/regTable[2][41] ) );
  LHQD1BWP \vrf/regTable_reg[2][42]  ( .E(n3589), .D(\vrf/N60 ), .Q(
        \vrf/regTable[2][42] ) );
  LHQD1BWP \vrf/regTable_reg[2][43]  ( .E(n3589), .D(\vrf/N61 ), .Q(
        \vrf/regTable[2][43] ) );
  LHQD1BWP \vrf/regTable_reg[2][44]  ( .E(n3589), .D(\vrf/N62 ), .Q(
        \vrf/regTable[2][44] ) );
  LHQD1BWP \vrf/regTable_reg[2][45]  ( .E(n3589), .D(\vrf/N63 ), .Q(
        \vrf/regTable[2][45] ) );
  LHQD1BWP \vrf/regTable_reg[2][46]  ( .E(n3589), .D(\vrf/N64 ), .Q(
        \vrf/regTable[2][46] ) );
  LHQD1BWP \vrf/regTable_reg[2][47]  ( .E(n3589), .D(\vrf/N65 ), .Q(
        \vrf/regTable[2][47] ) );
  LHQD1BWP \vrf/regTable_reg[2][48]  ( .E(n3589), .D(\vrf/N66 ), .Q(
        \vrf/regTable[2][48] ) );
  LHQD1BWP \vrf/regTable_reg[2][49]  ( .E(n3589), .D(\vrf/N67 ), .Q(
        \vrf/regTable[2][49] ) );
  LHQD1BWP \vrf/regTable_reg[2][50]  ( .E(n3589), .D(\vrf/N68 ), .Q(
        \vrf/regTable[2][50] ) );
  LHQD1BWP \vrf/regTable_reg[2][51]  ( .E(n3589), .D(\vrf/N69 ), .Q(
        \vrf/regTable[2][51] ) );
  LHQD1BWP \vrf/regTable_reg[2][52]  ( .E(n3589), .D(\vrf/N70 ), .Q(
        \vrf/regTable[2][52] ) );
  LHQD1BWP \vrf/regTable_reg[2][53]  ( .E(n3589), .D(\vrf/N71 ), .Q(
        \vrf/regTable[2][53] ) );
  LHQD1BWP \vrf/regTable_reg[2][54]  ( .E(n3589), .D(\vrf/N72 ), .Q(
        \vrf/regTable[2][54] ) );
  LHQD1BWP \vrf/regTable_reg[2][55]  ( .E(n3589), .D(\vrf/N73 ), .Q(
        \vrf/regTable[2][55] ) );
  LHQD1BWP \vrf/regTable_reg[2][56]  ( .E(n3589), .D(\vrf/N74 ), .Q(
        \vrf/regTable[2][56] ) );
  LHQD1BWP \vrf/regTable_reg[2][57]  ( .E(n3589), .D(\vrf/N75 ), .Q(
        \vrf/regTable[2][57] ) );
  LHQD1BWP \vrf/regTable_reg[2][58]  ( .E(n3589), .D(\vrf/N76 ), .Q(
        \vrf/regTable[2][58] ) );
  LHQD1BWP \vrf/regTable_reg[2][59]  ( .E(n3589), .D(\vrf/N77 ), .Q(
        \vrf/regTable[2][59] ) );
  LHQD1BWP \vrf/regTable_reg[2][60]  ( .E(n3589), .D(\vrf/N78 ), .Q(
        \vrf/regTable[2][60] ) );
  LHQD1BWP \vrf/regTable_reg[2][61]  ( .E(n3589), .D(\vrf/N79 ), .Q(
        \vrf/regTable[2][61] ) );
  LHQD1BWP \vrf/regTable_reg[2][62]  ( .E(n3589), .D(\vrf/N80 ), .Q(
        \vrf/regTable[2][62] ) );
  LHQD1BWP \vrf/regTable_reg[2][63]  ( .E(n3589), .D(\vrf/N81 ), .Q(
        \vrf/regTable[2][63] ) );
  LHQD1BWP \vrf/regTable_reg[2][64]  ( .E(n3589), .D(\vrf/N82 ), .Q(
        \vrf/regTable[2][64] ) );
  LHQD1BWP \vrf/regTable_reg[2][65]  ( .E(n3589), .D(\vrf/N83 ), .Q(
        \vrf/regTable[2][65] ) );
  LHQD1BWP \vrf/regTable_reg[2][66]  ( .E(n3589), .D(\vrf/N84 ), .Q(
        \vrf/regTable[2][66] ) );
  LHQD1BWP \vrf/regTable_reg[2][67]  ( .E(n3589), .D(\vrf/N85 ), .Q(
        \vrf/regTable[2][67] ) );
  LHQD1BWP \vrf/regTable_reg[2][68]  ( .E(n3589), .D(\vrf/N86 ), .Q(
        \vrf/regTable[2][68] ) );
  LHQD1BWP \vrf/regTable_reg[2][69]  ( .E(n3589), .D(\vrf/N87 ), .Q(
        \vrf/regTable[2][69] ) );
  LHQD1BWP \vrf/regTable_reg[2][70]  ( .E(n3589), .D(\vrf/N88 ), .Q(
        \vrf/regTable[2][70] ) );
  LHQD1BWP \vrf/regTable_reg[2][71]  ( .E(n3589), .D(\vrf/N89 ), .Q(
        \vrf/regTable[2][71] ) );
  LHQD1BWP \vrf/regTable_reg[2][72]  ( .E(n3589), .D(\vrf/N90 ), .Q(
        \vrf/regTable[2][72] ) );
  LHQD1BWP \vrf/regTable_reg[2][73]  ( .E(n3589), .D(\vrf/N91 ), .Q(
        \vrf/regTable[2][73] ) );
  LHQD1BWP \vrf/regTable_reg[2][74]  ( .E(n3589), .D(\vrf/N92 ), .Q(
        \vrf/regTable[2][74] ) );
  LHQD1BWP \vrf/regTable_reg[2][75]  ( .E(n3589), .D(\vrf/N93 ), .Q(
        \vrf/regTable[2][75] ) );
  LHQD1BWP \vrf/regTable_reg[2][76]  ( .E(n3589), .D(\vrf/N94 ), .Q(
        \vrf/regTable[2][76] ) );
  LHQD1BWP \vrf/regTable_reg[2][77]  ( .E(n3589), .D(\vrf/N95 ), .Q(
        \vrf/regTable[2][77] ) );
  LHQD1BWP \vrf/regTable_reg[2][78]  ( .E(n3589), .D(\vrf/N96 ), .Q(
        \vrf/regTable[2][78] ) );
  LHQD1BWP \vrf/regTable_reg[2][79]  ( .E(n3589), .D(\vrf/N97 ), .Q(
        \vrf/regTable[2][79] ) );
  LHQD1BWP \vrf/regTable_reg[2][80]  ( .E(n3589), .D(\vrf/N98 ), .Q(
        \vrf/regTable[2][80] ) );
  LHQD1BWP \vrf/regTable_reg[2][81]  ( .E(n3589), .D(\vrf/N99 ), .Q(
        \vrf/regTable[2][81] ) );
  LHQD1BWP \vrf/regTable_reg[2][82]  ( .E(n3589), .D(\vrf/N100 ), .Q(
        \vrf/regTable[2][82] ) );
  LHQD1BWP \vrf/regTable_reg[2][83]  ( .E(n3589), .D(\vrf/N101 ), .Q(
        \vrf/regTable[2][83] ) );
  LHQD1BWP \vrf/regTable_reg[2][84]  ( .E(n3589), .D(\vrf/N102 ), .Q(
        \vrf/regTable[2][84] ) );
  LHQD1BWP \vrf/regTable_reg[2][85]  ( .E(n3589), .D(\vrf/N103 ), .Q(
        \vrf/regTable[2][85] ) );
  LHQD1BWP \vrf/regTable_reg[2][86]  ( .E(n3589), .D(\vrf/N104 ), .Q(
        \vrf/regTable[2][86] ) );
  LHQD1BWP \vrf/regTable_reg[2][87]  ( .E(n3589), .D(\vrf/N105 ), .Q(
        \vrf/regTable[2][87] ) );
  LHQD1BWP \vrf/regTable_reg[2][88]  ( .E(n3589), .D(\vrf/N106 ), .Q(
        \vrf/regTable[2][88] ) );
  LHQD1BWP \vrf/regTable_reg[2][89]  ( .E(n3589), .D(\vrf/N107 ), .Q(
        \vrf/regTable[2][89] ) );
  LHQD1BWP \vrf/regTable_reg[2][90]  ( .E(n3589), .D(\vrf/N108 ), .Q(
        \vrf/regTable[2][90] ) );
  LHQD1BWP \vrf/regTable_reg[2][91]  ( .E(n3589), .D(\vrf/N109 ), .Q(
        \vrf/regTable[2][91] ) );
  LHQD1BWP \vrf/regTable_reg[2][92]  ( .E(n3589), .D(\vrf/N110 ), .Q(
        \vrf/regTable[2][92] ) );
  LHQD1BWP \vrf/regTable_reg[2][93]  ( .E(n3589), .D(\vrf/N111 ), .Q(
        \vrf/regTable[2][93] ) );
  LHQD1BWP \vrf/regTable_reg[2][94]  ( .E(n3589), .D(\vrf/N112 ), .Q(
        \vrf/regTable[2][94] ) );
  LHQD1BWP \vrf/regTable_reg[2][95]  ( .E(n3589), .D(\vrf/N113 ), .Q(
        \vrf/regTable[2][95] ) );
  LHQD1BWP \vrf/regTable_reg[2][96]  ( .E(n3589), .D(\vrf/N114 ), .Q(
        \vrf/regTable[2][96] ) );
  LHQD1BWP \vrf/regTable_reg[2][97]  ( .E(n3589), .D(\vrf/N115 ), .Q(
        \vrf/regTable[2][97] ) );
  LHQD1BWP \vrf/regTable_reg[2][98]  ( .E(n3589), .D(\vrf/N116 ), .Q(
        \vrf/regTable[2][98] ) );
  LHQD1BWP \vrf/regTable_reg[2][99]  ( .E(n3589), .D(\vrf/N118 ), .Q(
        \vrf/regTable[2][99] ) );
  LHQD1BWP \vrf/regTable_reg[2][100]  ( .E(n3589), .D(\vrf/N119 ), .Q(
        \vrf/regTable[2][100] ) );
  LHQD1BWP \vrf/regTable_reg[2][101]  ( .E(n3589), .D(\vrf/N120 ), .Q(
        \vrf/regTable[2][101] ) );
  LHQD1BWP \vrf/regTable_reg[2][102]  ( .E(n3589), .D(\vrf/N121 ), .Q(
        \vrf/regTable[2][102] ) );
  LHQD1BWP \vrf/regTable_reg[2][103]  ( .E(n3589), .D(\vrf/N122 ), .Q(
        \vrf/regTable[2][103] ) );
  LHQD1BWP \vrf/regTable_reg[2][104]  ( .E(n3589), .D(\vrf/N123 ), .Q(
        \vrf/regTable[2][104] ) );
  LHQD1BWP \vrf/regTable_reg[2][105]  ( .E(n3589), .D(\vrf/N124 ), .Q(
        \vrf/regTable[2][105] ) );
  LHQD1BWP \vrf/regTable_reg[2][106]  ( .E(n3589), .D(\vrf/N125 ), .Q(
        \vrf/regTable[2][106] ) );
  LHQD1BWP \vrf/regTable_reg[2][107]  ( .E(n3589), .D(\vrf/N126 ), .Q(
        \vrf/regTable[2][107] ) );
  LHQD1BWP \vrf/regTable_reg[2][108]  ( .E(n3589), .D(\vrf/N127 ), .Q(
        \vrf/regTable[2][108] ) );
  LHQD1BWP \vrf/regTable_reg[2][109]  ( .E(n3589), .D(\vrf/N128 ), .Q(
        \vrf/regTable[2][109] ) );
  LHQD1BWP \vrf/regTable_reg[2][110]  ( .E(n3589), .D(\vrf/N129 ), .Q(
        \vrf/regTable[2][110] ) );
  LHQD1BWP \vrf/regTable_reg[2][111]  ( .E(n3589), .D(\vrf/N130 ), .Q(
        \vrf/regTable[2][111] ) );
  LHQD1BWP \vrf/regTable_reg[2][112]  ( .E(n3589), .D(\vrf/N131 ), .Q(
        \vrf/regTable[2][112] ) );
  LHQD1BWP \vrf/regTable_reg[2][113]  ( .E(n3589), .D(\vrf/N132 ), .Q(
        \vrf/regTable[2][113] ) );
  LHQD1BWP \vrf/regTable_reg[2][114]  ( .E(n3589), .D(\vrf/N133 ), .Q(
        \vrf/regTable[2][114] ) );
  LHQD1BWP \vrf/regTable_reg[2][115]  ( .E(n3589), .D(\vrf/N134 ), .Q(
        \vrf/regTable[2][115] ) );
  LHQD1BWP \vrf/regTable_reg[2][116]  ( .E(n3589), .D(\vrf/N135 ), .Q(
        \vrf/regTable[2][116] ) );
  LHQD1BWP \vrf/regTable_reg[2][117]  ( .E(n3589), .D(\vrf/N136 ), .Q(
        \vrf/regTable[2][117] ) );
  LHQD1BWP \vrf/regTable_reg[2][118]  ( .E(n3589), .D(\vrf/N137 ), .Q(
        \vrf/regTable[2][118] ) );
  LHQD1BWP \vrf/regTable_reg[2][119]  ( .E(n3589), .D(\vrf/N138 ), .Q(
        \vrf/regTable[2][119] ) );
  LHQD1BWP \vrf/regTable_reg[2][120]  ( .E(n3589), .D(\vrf/N139 ), .Q(
        \vrf/regTable[2][120] ) );
  LHQD1BWP \vrf/regTable_reg[2][121]  ( .E(n3589), .D(\vrf/N140 ), .Q(
        \vrf/regTable[2][121] ) );
  LHQD1BWP \vrf/regTable_reg[2][122]  ( .E(n3589), .D(\vrf/N141 ), .Q(
        \vrf/regTable[2][122] ) );
  LHQD1BWP \vrf/regTable_reg[2][123]  ( .E(n3589), .D(\vrf/N142 ), .Q(
        \vrf/regTable[2][123] ) );
  LHQD1BWP \vrf/regTable_reg[2][124]  ( .E(n3589), .D(\vrf/N143 ), .Q(
        \vrf/regTable[2][124] ) );
  LHQD1BWP \vrf/regTable_reg[2][125]  ( .E(n3589), .D(\vrf/N144 ), .Q(
        \vrf/regTable[2][125] ) );
  LHQD1BWP \vrf/regTable_reg[2][126]  ( .E(n3589), .D(\vrf/N145 ), .Q(
        \vrf/regTable[2][126] ) );
  LHQD1BWP \vrf/regTable_reg[2][127]  ( .E(n3589), .D(\vrf/N146 ), .Q(
        \vrf/regTable[2][127] ) );
  LHQD1BWP \vrf/regTable_reg[2][128]  ( .E(n3589), .D(\vrf/N147 ), .Q(
        \vrf/regTable[2][128] ) );
  LHQD1BWP \vrf/regTable_reg[2][129]  ( .E(n3589), .D(\vrf/N148 ), .Q(
        \vrf/regTable[2][129] ) );
  LHQD1BWP \vrf/regTable_reg[2][130]  ( .E(n3589), .D(\vrf/N149 ), .Q(
        \vrf/regTable[2][130] ) );
  LHQD1BWP \vrf/regTable_reg[2][131]  ( .E(n3589), .D(\vrf/N150 ), .Q(
        \vrf/regTable[2][131] ) );
  LHQD1BWP \vrf/regTable_reg[2][132]  ( .E(n3589), .D(\vrf/N151 ), .Q(
        \vrf/regTable[2][132] ) );
  LHQD1BWP \vrf/regTable_reg[2][133]  ( .E(n3589), .D(\vrf/N152 ), .Q(
        \vrf/regTable[2][133] ) );
  LHQD1BWP \vrf/regTable_reg[2][134]  ( .E(n3589), .D(\vrf/N153 ), .Q(
        \vrf/regTable[2][134] ) );
  LHQD1BWP \vrf/regTable_reg[2][135]  ( .E(n3589), .D(\vrf/N154 ), .Q(
        \vrf/regTable[2][135] ) );
  LHQD1BWP \vrf/regTable_reg[2][136]  ( .E(n3589), .D(\vrf/N155 ), .Q(
        \vrf/regTable[2][136] ) );
  LHQD1BWP \vrf/regTable_reg[2][137]  ( .E(\vrf/N290 ), .D(\vrf/N156 ), .Q(
        \vrf/regTable[2][137] ) );
  LHQD1BWP \vrf/regTable_reg[2][138]  ( .E(n3589), .D(\vrf/N157 ), .Q(
        \vrf/regTable[2][138] ) );
  LHQD1BWP \vrf/regTable_reg[2][139]  ( .E(\vrf/N290 ), .D(\vrf/N158 ), .Q(
        \vrf/regTable[2][139] ) );
  LHQD1BWP \vrf/regTable_reg[2][140]  ( .E(n3589), .D(\vrf/N159 ), .Q(
        \vrf/regTable[2][140] ) );
  LHQD1BWP \vrf/regTable_reg[2][141]  ( .E(\vrf/N290 ), .D(\vrf/N160 ), .Q(
        \vrf/regTable[2][141] ) );
  LHQD1BWP \vrf/regTable_reg[2][142]  ( .E(n3589), .D(\vrf/N161 ), .Q(
        \vrf/regTable[2][142] ) );
  LHQD1BWP \vrf/regTable_reg[2][143]  ( .E(\vrf/N290 ), .D(\vrf/N162 ), .Q(
        \vrf/regTable[2][143] ) );
  LHQD1BWP \vrf/regTable_reg[2][144]  ( .E(n3589), .D(\vrf/N163 ), .Q(
        \vrf/regTable[2][144] ) );
  LHQD1BWP \vrf/regTable_reg[2][145]  ( .E(\vrf/N290 ), .D(\vrf/N164 ), .Q(
        \vrf/regTable[2][145] ) );
  LHQD1BWP \vrf/regTable_reg[2][146]  ( .E(n3589), .D(\vrf/N165 ), .Q(
        \vrf/regTable[2][146] ) );
  LHQD1BWP \vrf/regTable_reg[2][147]  ( .E(\vrf/N290 ), .D(\vrf/N166 ), .Q(
        \vrf/regTable[2][147] ) );
  LHQD1BWP \vrf/regTable_reg[2][148]  ( .E(n3589), .D(\vrf/N167 ), .Q(
        \vrf/regTable[2][148] ) );
  LHQD1BWP \vrf/regTable_reg[2][149]  ( .E(n3589), .D(\vrf/N168 ), .Q(
        \vrf/regTable[2][149] ) );
  LHQD1BWP \vrf/regTable_reg[2][150]  ( .E(n3589), .D(\vrf/N169 ), .Q(
        \vrf/regTable[2][150] ) );
  LHQD1BWP \vrf/regTable_reg[2][151]  ( .E(\vrf/N290 ), .D(\vrf/N170 ), .Q(
        \vrf/regTable[2][151] ) );
  LHQD1BWP \vrf/regTable_reg[2][152]  ( .E(n3589), .D(\vrf/N171 ), .Q(
        \vrf/regTable[2][152] ) );
  LHQD1BWP \vrf/regTable_reg[2][153]  ( .E(n3589), .D(\vrf/N172 ), .Q(
        \vrf/regTable[2][153] ) );
  LHQD1BWP \vrf/regTable_reg[2][154]  ( .E(n3589), .D(\vrf/N173 ), .Q(
        \vrf/regTable[2][154] ) );
  LHQD1BWP \vrf/regTable_reg[2][155]  ( .E(\vrf/N290 ), .D(\vrf/N174 ), .Q(
        \vrf/regTable[2][155] ) );
  LHQD1BWP \vrf/regTable_reg[2][156]  ( .E(n3589), .D(\vrf/N175 ), .Q(
        \vrf/regTable[2][156] ) );
  LHQD1BWP \vrf/regTable_reg[2][157]  ( .E(n3589), .D(\vrf/N176 ), .Q(
        \vrf/regTable[2][157] ) );
  LHQD1BWP \vrf/regTable_reg[2][158]  ( .E(n3589), .D(\vrf/N177 ), .Q(
        \vrf/regTable[2][158] ) );
  LHQD1BWP \vrf/regTable_reg[2][159]  ( .E(n3589), .D(\vrf/N178 ), .Q(
        \vrf/regTable[2][159] ) );
  LHQD1BWP \vrf/regTable_reg[2][160]  ( .E(\vrf/N290 ), .D(\vrf/N179 ), .Q(
        \vrf/regTable[2][160] ) );
  LHQD1BWP \vrf/regTable_reg[2][161]  ( .E(n3589), .D(\vrf/N180 ), .Q(
        \vrf/regTable[2][161] ) );
  LHQD1BWP \vrf/regTable_reg[2][162]  ( .E(n3589), .D(\vrf/N181 ), .Q(
        \vrf/regTable[2][162] ) );
  LHQD1BWP \vrf/regTable_reg[2][163]  ( .E(n3589), .D(\vrf/N182 ), .Q(
        \vrf/regTable[2][163] ) );
  LHQD1BWP \vrf/regTable_reg[2][164]  ( .E(\vrf/N290 ), .D(\vrf/N183 ), .Q(
        \vrf/regTable[2][164] ) );
  LHQD1BWP \vrf/regTable_reg[2][165]  ( .E(n3589), .D(\vrf/N184 ), .Q(
        \vrf/regTable[2][165] ) );
  LHQD1BWP \vrf/regTable_reg[2][166]  ( .E(n3589), .D(\vrf/N185 ), .Q(
        \vrf/regTable[2][166] ) );
  LHQD1BWP \vrf/regTable_reg[2][167]  ( .E(n3589), .D(\vrf/N186 ), .Q(
        \vrf/regTable[2][167] ) );
  LHQD1BWP \vrf/regTable_reg[2][168]  ( .E(\vrf/N290 ), .D(\vrf/N187 ), .Q(
        \vrf/regTable[2][168] ) );
  LHQD1BWP \vrf/regTable_reg[2][169]  ( .E(n3589), .D(\vrf/N188 ), .Q(
        \vrf/regTable[2][169] ) );
  LHQD1BWP \vrf/regTable_reg[2][170]  ( .E(n3589), .D(\vrf/N189 ), .Q(
        \vrf/regTable[2][170] ) );
  LHQD1BWP \vrf/regTable_reg[2][171]  ( .E(n3589), .D(\vrf/N190 ), .Q(
        \vrf/regTable[2][171] ) );
  LHQD1BWP \vrf/regTable_reg[2][172]  ( .E(n3589), .D(\vrf/N191 ), .Q(
        \vrf/regTable[2][172] ) );
  LHQD1BWP \vrf/regTable_reg[2][173]  ( .E(n3589), .D(\vrf/N192 ), .Q(
        \vrf/regTable[2][173] ) );
  LHQD1BWP \vrf/regTable_reg[2][174]  ( .E(\vrf/N290 ), .D(\vrf/N193 ), .Q(
        \vrf/regTable[2][174] ) );
  LHQD1BWP \vrf/regTable_reg[2][175]  ( .E(n3589), .D(\vrf/N194 ), .Q(
        \vrf/regTable[2][175] ) );
  LHQD1BWP \vrf/regTable_reg[2][176]  ( .E(n3589), .D(\vrf/N195 ), .Q(
        \vrf/regTable[2][176] ) );
  LHQD1BWP \vrf/regTable_reg[2][177]  ( .E(n3589), .D(\vrf/N196 ), .Q(
        \vrf/regTable[2][177] ) );
  LHQD1BWP \vrf/regTable_reg[2][178]  ( .E(n3589), .D(\vrf/N197 ), .Q(
        \vrf/regTable[2][178] ) );
  LHQD1BWP \vrf/regTable_reg[2][179]  ( .E(\vrf/N290 ), .D(\vrf/N198 ), .Q(
        \vrf/regTable[2][179] ) );
  LHQD1BWP \vrf/regTable_reg[2][180]  ( .E(n3589), .D(\vrf/N199 ), .Q(
        \vrf/regTable[2][180] ) );
  LHQD1BWP \vrf/regTable_reg[2][181]  ( .E(n3589), .D(\vrf/N200 ), .Q(
        \vrf/regTable[2][181] ) );
  LHQD1BWP \vrf/regTable_reg[2][182]  ( .E(n3589), .D(\vrf/N201 ), .Q(
        \vrf/regTable[2][182] ) );
  LHQD1BWP \vrf/regTable_reg[2][183]  ( .E(n3589), .D(\vrf/N202 ), .Q(
        \vrf/regTable[2][183] ) );
  LHQD1BWP \vrf/regTable_reg[2][184]  ( .E(n3589), .D(\vrf/N203 ), .Q(
        \vrf/regTable[2][184] ) );
  LHQD1BWP \vrf/regTable_reg[2][185]  ( .E(n3589), .D(\vrf/N204 ), .Q(
        \vrf/regTable[2][185] ) );
  LHQD1BWP \vrf/regTable_reg[2][186]  ( .E(n3589), .D(\vrf/N205 ), .Q(
        \vrf/regTable[2][186] ) );
  LHQD1BWP \vrf/regTable_reg[2][187]  ( .E(n3589), .D(\vrf/N206 ), .Q(
        \vrf/regTable[2][187] ) );
  LHQD1BWP \vrf/regTable_reg[2][188]  ( .E(n3589), .D(\vrf/N207 ), .Q(
        \vrf/regTable[2][188] ) );
  LHQD1BWP \vrf/regTable_reg[2][189]  ( .E(\vrf/N290 ), .D(\vrf/N208 ), .Q(
        \vrf/regTable[2][189] ) );
  LHQD1BWP \vrf/regTable_reg[2][190]  ( .E(n3589), .D(\vrf/N209 ), .Q(
        \vrf/regTable[2][190] ) );
  LHQD1BWP \vrf/regTable_reg[2][191]  ( .E(n3589), .D(\vrf/N210 ), .Q(
        \vrf/regTable[2][191] ) );
  LHQD1BWP \vrf/regTable_reg[2][192]  ( .E(n3589), .D(\vrf/N211 ), .Q(
        \vrf/regTable[2][192] ) );
  LHQD1BWP \vrf/regTable_reg[2][193]  ( .E(n3589), .D(\vrf/N212 ), .Q(
        \vrf/regTable[2][193] ) );
  LHQD1BWP \vrf/regTable_reg[2][194]  ( .E(\vrf/N290 ), .D(\vrf/N213 ), .Q(
        \vrf/regTable[2][194] ) );
  LHQD1BWP \vrf/regTable_reg[2][195]  ( .E(\vrf/N290 ), .D(\vrf/N214 ), .Q(
        \vrf/regTable[2][195] ) );
  LHQD1BWP \vrf/regTable_reg[2][196]  ( .E(n3589), .D(\vrf/N215 ), .Q(
        \vrf/regTable[2][196] ) );
  LHQD1BWP \vrf/regTable_reg[2][197]  ( .E(n3589), .D(\vrf/N216 ), .Q(
        \vrf/regTable[2][197] ) );
  LHQD1BWP \vrf/regTable_reg[2][198]  ( .E(n3589), .D(\vrf/N218 ), .Q(
        \vrf/regTable[2][198] ) );
  LHQD1BWP \vrf/regTable_reg[2][199]  ( .E(n3589), .D(\vrf/N219 ), .Q(
        \vrf/regTable[2][199] ) );
  LHQD1BWP \vrf/regTable_reg[2][200]  ( .E(n3589), .D(\vrf/N220 ), .Q(
        \vrf/regTable[2][200] ) );
  LHQD1BWP \vrf/regTable_reg[2][201]  ( .E(\vrf/N290 ), .D(\vrf/N221 ), .Q(
        \vrf/regTable[2][201] ) );
  LHQD1BWP \vrf/regTable_reg[2][202]  ( .E(n3589), .D(\vrf/N222 ), .Q(
        \vrf/regTable[2][202] ) );
  LHQD1BWP \vrf/regTable_reg[2][203]  ( .E(n3589), .D(\vrf/N223 ), .Q(
        \vrf/regTable[2][203] ) );
  LHQD1BWP \vrf/regTable_reg[2][204]  ( .E(\vrf/N290 ), .D(\vrf/N224 ), .Q(
        \vrf/regTable[2][204] ) );
  LHQD1BWP \vrf/regTable_reg[2][205]  ( .E(n3589), .D(\vrf/N225 ), .Q(
        \vrf/regTable[2][205] ) );
  LHQD1BWP \vrf/regTable_reg[2][206]  ( .E(\vrf/N290 ), .D(\vrf/N226 ), .Q(
        \vrf/regTable[2][206] ) );
  LHQD1BWP \vrf/regTable_reg[2][207]  ( .E(n3589), .D(\vrf/N227 ), .Q(
        \vrf/regTable[2][207] ) );
  LHQD1BWP \vrf/regTable_reg[2][208]  ( .E(n3589), .D(\vrf/N228 ), .Q(
        \vrf/regTable[2][208] ) );
  LHQD1BWP \vrf/regTable_reg[2][209]  ( .E(n3589), .D(\vrf/N229 ), .Q(
        \vrf/regTable[2][209] ) );
  LHQD1BWP \vrf/regTable_reg[2][210]  ( .E(n3589), .D(\vrf/N230 ), .Q(
        \vrf/regTable[2][210] ) );
  LHQD1BWP \vrf/regTable_reg[2][211]  ( .E(n3589), .D(\vrf/N231 ), .Q(
        \vrf/regTable[2][211] ) );
  LHQD1BWP \vrf/regTable_reg[2][212]  ( .E(n3589), .D(\vrf/N232 ), .Q(
        \vrf/regTable[2][212] ) );
  LHQD1BWP \vrf/regTable_reg[2][213]  ( .E(n3589), .D(\vrf/N233 ), .Q(
        \vrf/regTable[2][213] ) );
  LHQD1BWP \vrf/regTable_reg[2][214]  ( .E(n3589), .D(\vrf/N234 ), .Q(
        \vrf/regTable[2][214] ) );
  LHQD1BWP \vrf/regTable_reg[2][215]  ( .E(n3589), .D(\vrf/N235 ), .Q(
        \vrf/regTable[2][215] ) );
  LHQD1BWP \vrf/regTable_reg[2][216]  ( .E(n3589), .D(\vrf/N236 ), .Q(
        \vrf/regTable[2][216] ) );
  LHQD1BWP \vrf/regTable_reg[2][217]  ( .E(n3589), .D(\vrf/N237 ), .Q(
        \vrf/regTable[2][217] ) );
  LHQD1BWP \vrf/regTable_reg[2][218]  ( .E(n3589), .D(\vrf/N238 ), .Q(
        \vrf/regTable[2][218] ) );
  LHQD1BWP \vrf/regTable_reg[2][219]  ( .E(n3589), .D(\vrf/N239 ), .Q(
        \vrf/regTable[2][219] ) );
  LHQD1BWP \vrf/regTable_reg[2][220]  ( .E(n3589), .D(\vrf/N240 ), .Q(
        \vrf/regTable[2][220] ) );
  LHQD1BWP \vrf/regTable_reg[2][221]  ( .E(n3589), .D(\vrf/N241 ), .Q(
        \vrf/regTable[2][221] ) );
  LHQD1BWP \vrf/regTable_reg[2][222]  ( .E(n3589), .D(\vrf/N242 ), .Q(
        \vrf/regTable[2][222] ) );
  LHQD1BWP \vrf/regTable_reg[2][223]  ( .E(\vrf/N290 ), .D(\vrf/N243 ), .Q(
        \vrf/regTable[2][223] ) );
  LHQD1BWP \vrf/regTable_reg[2][224]  ( .E(n3589), .D(\vrf/N244 ), .Q(
        \vrf/regTable[2][224] ) );
  LHQD1BWP \vrf/regTable_reg[2][225]  ( .E(n3589), .D(\vrf/N245 ), .Q(
        \vrf/regTable[2][225] ) );
  LHQD1BWP \vrf/regTable_reg[2][226]  ( .E(n3589), .D(\vrf/N246 ), .Q(
        \vrf/regTable[2][226] ) );
  LHQD1BWP \vrf/regTable_reg[2][227]  ( .E(\vrf/N290 ), .D(\vrf/N247 ), .Q(
        \vrf/regTable[2][227] ) );
  LHQD1BWP \vrf/regTable_reg[2][228]  ( .E(n3589), .D(\vrf/N248 ), .Q(
        \vrf/regTable[2][228] ) );
  LHQD1BWP \vrf/regTable_reg[2][229]  ( .E(n3589), .D(\vrf/N249 ), .Q(
        \vrf/regTable[2][229] ) );
  LHQD1BWP \vrf/regTable_reg[2][230]  ( .E(n3589), .D(\vrf/N250 ), .Q(
        \vrf/regTable[2][230] ) );
  LHQD1BWP \vrf/regTable_reg[2][231]  ( .E(\vrf/N290 ), .D(\vrf/N251 ), .Q(
        \vrf/regTable[2][231] ) );
  LHQD1BWP \vrf/regTable_reg[2][232]  ( .E(n3589), .D(\vrf/N252 ), .Q(
        \vrf/regTable[2][232] ) );
  LHQD1BWP \vrf/regTable_reg[2][233]  ( .E(n3589), .D(\vrf/N253 ), .Q(
        \vrf/regTable[2][233] ) );
  LHQD1BWP \vrf/regTable_reg[2][234]  ( .E(n3589), .D(\vrf/N254 ), .Q(
        \vrf/regTable[2][234] ) );
  LHQD1BWP \vrf/regTable_reg[2][235]  ( .E(n3589), .D(\vrf/N255 ), .Q(
        \vrf/regTable[2][235] ) );
  LHQD1BWP \vrf/regTable_reg[2][236]  ( .E(n3589), .D(\vrf/N256 ), .Q(
        \vrf/regTable[2][236] ) );
  LHQD1BWP \vrf/regTable_reg[2][237]  ( .E(n3589), .D(\vrf/N257 ), .Q(
        \vrf/regTable[2][237] ) );
  LHQD1BWP \vrf/regTable_reg[2][238]  ( .E(n3589), .D(\vrf/N258 ), .Q(
        \vrf/regTable[2][238] ) );
  LHQD1BWP \vrf/regTable_reg[2][239]  ( .E(n3589), .D(\vrf/N259 ), .Q(
        \vrf/regTable[2][239] ) );
  LHQD1BWP \vrf/regTable_reg[2][240]  ( .E(n3589), .D(\vrf/N260 ), .Q(
        \vrf/regTable[2][240] ) );
  LHQD1BWP \vrf/regTable_reg[2][241]  ( .E(n3589), .D(\vrf/N261 ), .Q(
        \vrf/regTable[2][241] ) );
  LHQD1BWP \vrf/regTable_reg[2][242]  ( .E(n3589), .D(\vrf/N262 ), .Q(
        \vrf/regTable[2][242] ) );
  LHQD1BWP \vrf/regTable_reg[2][243]  ( .E(n3589), .D(\vrf/N263 ), .Q(
        \vrf/regTable[2][243] ) );
  LHQD1BWP \vrf/regTable_reg[2][244]  ( .E(n3589), .D(\vrf/N264 ), .Q(
        \vrf/regTable[2][244] ) );
  LHQD1BWP \vrf/regTable_reg[2][245]  ( .E(n3589), .D(\vrf/N265 ), .Q(
        \vrf/regTable[2][245] ) );
  LHQD1BWP \vrf/regTable_reg[2][246]  ( .E(n3589), .D(\vrf/N266 ), .Q(
        \vrf/regTable[2][246] ) );
  LHQD1BWP \vrf/regTable_reg[2][247]  ( .E(n3589), .D(\vrf/N267 ), .Q(
        \vrf/regTable[2][247] ) );
  LHQD1BWP \vrf/regTable_reg[2][248]  ( .E(n3589), .D(\vrf/N268 ), .Q(
        \vrf/regTable[2][248] ) );
  LHQD1BWP \vrf/regTable_reg[2][249]  ( .E(n3589), .D(\vrf/N269 ), .Q(
        \vrf/regTable[2][249] ) );
  LHQD1BWP \vrf/regTable_reg[2][250]  ( .E(n3589), .D(\vrf/N270 ), .Q(
        \vrf/regTable[2][250] ) );
  LHQD1BWP \vrf/regTable_reg[2][251]  ( .E(\vrf/N290 ), .D(\vrf/N271 ), .Q(
        \vrf/regTable[2][251] ) );
  LHQD1BWP \vrf/regTable_reg[2][252]  ( .E(n3589), .D(\vrf/N272 ), .Q(
        \vrf/regTable[2][252] ) );
  LHQD1BWP \vrf/regTable_reg[2][253]  ( .E(n3589), .D(\vrf/N273 ), .Q(
        \vrf/regTable[2][253] ) );
  LHQD1BWP \vrf/regTable_reg[2][254]  ( .E(n3589), .D(\vrf/N274 ), .Q(
        \vrf/regTable[2][254] ) );
  LHQD1BWP \vrf/regTable_reg[2][255]  ( .E(n3589), .D(\vrf/N275 ), .Q(
        \vrf/regTable[2][255] ) );
  LHQD1BWP \vrf/regTable_reg[1][0]  ( .E(n3588), .D(\vrf/N18 ), .Q(
        \vrf/regTable[1][0] ) );
  LHQD1BWP \vrf/regTable_reg[1][1]  ( .E(n3588), .D(\vrf/N19 ), .Q(
        \vrf/regTable[1][1] ) );
  LHQD1BWP \vrf/regTable_reg[1][2]  ( .E(n3588), .D(\vrf/N20 ), .Q(
        \vrf/regTable[1][2] ) );
  LHQD1BWP \vrf/regTable_reg[1][3]  ( .E(n3588), .D(\vrf/N21 ), .Q(
        \vrf/regTable[1][3] ) );
  LHQD1BWP \vrf/regTable_reg[1][4]  ( .E(n3588), .D(\vrf/N22 ), .Q(
        \vrf/regTable[1][4] ) );
  LHQD1BWP \vrf/regTable_reg[1][5]  ( .E(n3588), .D(\vrf/N23 ), .Q(
        \vrf/regTable[1][5] ) );
  LHQD1BWP \vrf/regTable_reg[1][6]  ( .E(n3588), .D(\vrf/N24 ), .Q(
        \vrf/regTable[1][6] ) );
  LHQD1BWP \vrf/regTable_reg[1][7]  ( .E(n3588), .D(\vrf/N25 ), .Q(
        \vrf/regTable[1][7] ) );
  LHQD1BWP \vrf/regTable_reg[1][8]  ( .E(n3588), .D(\vrf/N26 ), .Q(
        \vrf/regTable[1][8] ) );
  LHQD1BWP \vrf/regTable_reg[1][9]  ( .E(n3588), .D(\vrf/N27 ), .Q(
        \vrf/regTable[1][9] ) );
  LHQD1BWP \vrf/regTable_reg[1][10]  ( .E(n3588), .D(\vrf/N28 ), .Q(
        \vrf/regTable[1][10] ) );
  LHQD1BWP \vrf/regTable_reg[1][11]  ( .E(n3588), .D(\vrf/N29 ), .Q(
        \vrf/regTable[1][11] ) );
  LHQD1BWP \vrf/regTable_reg[1][12]  ( .E(n3588), .D(\vrf/N30 ), .Q(
        \vrf/regTable[1][12] ) );
  LHQD1BWP \vrf/regTable_reg[1][13]  ( .E(n3588), .D(\vrf/N31 ), .Q(
        \vrf/regTable[1][13] ) );
  LHQD1BWP \vrf/regTable_reg[1][14]  ( .E(n3588), .D(\vrf/N32 ), .Q(
        \vrf/regTable[1][14] ) );
  LHQD1BWP \vrf/regTable_reg[1][15]  ( .E(n3588), .D(\vrf/N33 ), .Q(
        \vrf/regTable[1][15] ) );
  LHQD1BWP \vrf/regTable_reg[1][16]  ( .E(n3588), .D(\vrf/N34 ), .Q(
        \vrf/regTable[1][16] ) );
  LHQD1BWP \vrf/regTable_reg[1][17]  ( .E(n3588), .D(\vrf/N35 ), .Q(
        \vrf/regTable[1][17] ) );
  LHQD1BWP \vrf/regTable_reg[1][18]  ( .E(n3588), .D(\vrf/N36 ), .Q(
        \vrf/regTable[1][18] ) );
  LHQD1BWP \vrf/regTable_reg[1][19]  ( .E(n3588), .D(\vrf/N37 ), .Q(
        \vrf/regTable[1][19] ) );
  LHQD1BWP \vrf/regTable_reg[1][20]  ( .E(n3588), .D(\vrf/N38 ), .Q(
        \vrf/regTable[1][20] ) );
  LHQD1BWP \vrf/regTable_reg[1][21]  ( .E(n3588), .D(\vrf/N39 ), .Q(
        \vrf/regTable[1][21] ) );
  LHQD1BWP \vrf/regTable_reg[1][22]  ( .E(n3588), .D(\vrf/N40 ), .Q(
        \vrf/regTable[1][22] ) );
  LHQD1BWP \vrf/regTable_reg[1][23]  ( .E(n3588), .D(\vrf/N41 ), .Q(
        \vrf/regTable[1][23] ) );
  LHQD1BWP \vrf/regTable_reg[1][24]  ( .E(n3588), .D(\vrf/N42 ), .Q(
        \vrf/regTable[1][24] ) );
  LHQD1BWP \vrf/regTable_reg[1][25]  ( .E(n3588), .D(\vrf/N43 ), .Q(
        \vrf/regTable[1][25] ) );
  LHQD1BWP \vrf/regTable_reg[1][26]  ( .E(n3588), .D(\vrf/N44 ), .Q(
        \vrf/regTable[1][26] ) );
  LHQD1BWP \vrf/regTable_reg[1][27]  ( .E(n3588), .D(\vrf/N45 ), .Q(
        \vrf/regTable[1][27] ) );
  LHQD1BWP \vrf/regTable_reg[1][28]  ( .E(n3588), .D(\vrf/N46 ), .Q(
        \vrf/regTable[1][28] ) );
  LHQD1BWP \vrf/regTable_reg[1][29]  ( .E(n3588), .D(\vrf/N47 ), .Q(
        \vrf/regTable[1][29] ) );
  LHQD1BWP \vrf/regTable_reg[1][30]  ( .E(n3588), .D(\vrf/N48 ), .Q(
        \vrf/regTable[1][30] ) );
  LHQD1BWP \vrf/regTable_reg[1][31]  ( .E(n3588), .D(\vrf/N49 ), .Q(
        \vrf/regTable[1][31] ) );
  LHQD1BWP \vrf/regTable_reg[1][32]  ( .E(n3588), .D(\vrf/N50 ), .Q(
        \vrf/regTable[1][32] ) );
  LHQD1BWP \vrf/regTable_reg[1][33]  ( .E(n3588), .D(\vrf/N51 ), .Q(
        \vrf/regTable[1][33] ) );
  LHQD1BWP \vrf/regTable_reg[1][34]  ( .E(n3588), .D(\vrf/N52 ), .Q(
        \vrf/regTable[1][34] ) );
  LHQD1BWP \vrf/regTable_reg[1][35]  ( .E(n3588), .D(\vrf/N53 ), .Q(
        \vrf/regTable[1][35] ) );
  LHQD1BWP \vrf/regTable_reg[1][36]  ( .E(n3588), .D(\vrf/N54 ), .Q(
        \vrf/regTable[1][36] ) );
  LHQD1BWP \vrf/regTable_reg[1][37]  ( .E(n3588), .D(\vrf/N55 ), .Q(
        \vrf/regTable[1][37] ) );
  LHQD1BWP \vrf/regTable_reg[1][38]  ( .E(n3588), .D(\vrf/N56 ), .Q(
        \vrf/regTable[1][38] ) );
  LHQD1BWP \vrf/regTable_reg[1][39]  ( .E(n3588), .D(\vrf/N57 ), .Q(
        \vrf/regTable[1][39] ) );
  LHQD1BWP \vrf/regTable_reg[1][40]  ( .E(n3588), .D(\vrf/N58 ), .Q(
        \vrf/regTable[1][40] ) );
  LHQD1BWP \vrf/regTable_reg[1][41]  ( .E(n3588), .D(\vrf/N59 ), .Q(
        \vrf/regTable[1][41] ) );
  LHQD1BWP \vrf/regTable_reg[1][42]  ( .E(n3588), .D(\vrf/N60 ), .Q(
        \vrf/regTable[1][42] ) );
  LHQD1BWP \vrf/regTable_reg[1][43]  ( .E(n3588), .D(\vrf/N61 ), .Q(
        \vrf/regTable[1][43] ) );
  LHQD1BWP \vrf/regTable_reg[1][44]  ( .E(n3588), .D(\vrf/N62 ), .Q(
        \vrf/regTable[1][44] ) );
  LHQD1BWP \vrf/regTable_reg[1][45]  ( .E(n3588), .D(\vrf/N63 ), .Q(
        \vrf/regTable[1][45] ) );
  LHQD1BWP \vrf/regTable_reg[1][46]  ( .E(n3588), .D(\vrf/N64 ), .Q(
        \vrf/regTable[1][46] ) );
  LHQD1BWP \vrf/regTable_reg[1][47]  ( .E(n3588), .D(\vrf/N65 ), .Q(
        \vrf/regTable[1][47] ) );
  LHQD1BWP \vrf/regTable_reg[1][48]  ( .E(n3588), .D(\vrf/N66 ), .Q(
        \vrf/regTable[1][48] ) );
  LHQD1BWP \vrf/regTable_reg[1][49]  ( .E(n3588), .D(\vrf/N67 ), .Q(
        \vrf/regTable[1][49] ) );
  LHQD1BWP \vrf/regTable_reg[1][50]  ( .E(n3588), .D(\vrf/N68 ), .Q(
        \vrf/regTable[1][50] ) );
  LHQD1BWP \vrf/regTable_reg[1][51]  ( .E(n3588), .D(\vrf/N69 ), .Q(
        \vrf/regTable[1][51] ) );
  LHQD1BWP \vrf/regTable_reg[1][52]  ( .E(n3588), .D(\vrf/N70 ), .Q(
        \vrf/regTable[1][52] ) );
  LHQD1BWP \vrf/regTable_reg[1][53]  ( .E(n3588), .D(\vrf/N71 ), .Q(
        \vrf/regTable[1][53] ) );
  LHQD1BWP \vrf/regTable_reg[1][54]  ( .E(n3588), .D(\vrf/N72 ), .Q(
        \vrf/regTable[1][54] ) );
  LHQD1BWP \vrf/regTable_reg[1][55]  ( .E(n3588), .D(\vrf/N73 ), .Q(
        \vrf/regTable[1][55] ) );
  LHQD1BWP \vrf/regTable_reg[1][56]  ( .E(n3588), .D(\vrf/N74 ), .Q(
        \vrf/regTable[1][56] ) );
  LHQD1BWP \vrf/regTable_reg[1][57]  ( .E(n3588), .D(\vrf/N75 ), .Q(
        \vrf/regTable[1][57] ) );
  LHQD1BWP \vrf/regTable_reg[1][58]  ( .E(n3588), .D(\vrf/N76 ), .Q(
        \vrf/regTable[1][58] ) );
  LHQD1BWP \vrf/regTable_reg[1][59]  ( .E(n3588), .D(\vrf/N77 ), .Q(
        \vrf/regTable[1][59] ) );
  LHQD1BWP \vrf/regTable_reg[1][60]  ( .E(n3588), .D(\vrf/N78 ), .Q(
        \vrf/regTable[1][60] ) );
  LHQD1BWP \vrf/regTable_reg[1][61]  ( .E(n3588), .D(\vrf/N79 ), .Q(
        \vrf/regTable[1][61] ) );
  LHQD1BWP \vrf/regTable_reg[1][62]  ( .E(n3588), .D(\vrf/N80 ), .Q(
        \vrf/regTable[1][62] ) );
  LHQD1BWP \vrf/regTable_reg[1][63]  ( .E(n3588), .D(\vrf/N81 ), .Q(
        \vrf/regTable[1][63] ) );
  LHQD1BWP \vrf/regTable_reg[1][64]  ( .E(n3588), .D(\vrf/N82 ), .Q(
        \vrf/regTable[1][64] ) );
  LHQD1BWP \vrf/regTable_reg[1][65]  ( .E(n3588), .D(\vrf/N83 ), .Q(
        \vrf/regTable[1][65] ) );
  LHQD1BWP \vrf/regTable_reg[1][66]  ( .E(n3588), .D(\vrf/N84 ), .Q(
        \vrf/regTable[1][66] ) );
  LHQD1BWP \vrf/regTable_reg[1][67]  ( .E(n3588), .D(\vrf/N85 ), .Q(
        \vrf/regTable[1][67] ) );
  LHQD1BWP \vrf/regTable_reg[1][68]  ( .E(n3588), .D(\vrf/N86 ), .Q(
        \vrf/regTable[1][68] ) );
  LHQD1BWP \vrf/regTable_reg[1][69]  ( .E(n3588), .D(\vrf/N87 ), .Q(
        \vrf/regTable[1][69] ) );
  LHQD1BWP \vrf/regTable_reg[1][70]  ( .E(n3588), .D(\vrf/N88 ), .Q(
        \vrf/regTable[1][70] ) );
  LHQD1BWP \vrf/regTable_reg[1][71]  ( .E(n3588), .D(\vrf/N89 ), .Q(
        \vrf/regTable[1][71] ) );
  LHQD1BWP \vrf/regTable_reg[1][72]  ( .E(n3588), .D(\vrf/N90 ), .Q(
        \vrf/regTable[1][72] ) );
  LHQD1BWP \vrf/regTable_reg[1][73]  ( .E(n3588), .D(\vrf/N91 ), .Q(
        \vrf/regTable[1][73] ) );
  LHQD1BWP \vrf/regTable_reg[1][74]  ( .E(n3588), .D(\vrf/N92 ), .Q(
        \vrf/regTable[1][74] ) );
  LHQD1BWP \vrf/regTable_reg[1][75]  ( .E(n3588), .D(\vrf/N93 ), .Q(
        \vrf/regTable[1][75] ) );
  LHQD1BWP \vrf/regTable_reg[1][76]  ( .E(n3588), .D(\vrf/N94 ), .Q(
        \vrf/regTable[1][76] ) );
  LHQD1BWP \vrf/regTable_reg[1][77]  ( .E(n3588), .D(\vrf/N95 ), .Q(
        \vrf/regTable[1][77] ) );
  LHQD1BWP \vrf/regTable_reg[1][78]  ( .E(n3588), .D(\vrf/N96 ), .Q(
        \vrf/regTable[1][78] ) );
  LHQD1BWP \vrf/regTable_reg[1][79]  ( .E(n3588), .D(\vrf/N97 ), .Q(
        \vrf/regTable[1][79] ) );
  LHQD1BWP \vrf/regTable_reg[1][80]  ( .E(n3588), .D(\vrf/N98 ), .Q(
        \vrf/regTable[1][80] ) );
  LHQD1BWP \vrf/regTable_reg[1][81]  ( .E(n3588), .D(\vrf/N99 ), .Q(
        \vrf/regTable[1][81] ) );
  LHQD1BWP \vrf/regTable_reg[1][82]  ( .E(n3588), .D(\vrf/N100 ), .Q(
        \vrf/regTable[1][82] ) );
  LHQD1BWP \vrf/regTable_reg[1][83]  ( .E(n3588), .D(\vrf/N101 ), .Q(
        \vrf/regTable[1][83] ) );
  LHQD1BWP \vrf/regTable_reg[1][84]  ( .E(n3588), .D(\vrf/N102 ), .Q(
        \vrf/regTable[1][84] ) );
  LHQD1BWP \vrf/regTable_reg[1][85]  ( .E(n3588), .D(\vrf/N103 ), .Q(
        \vrf/regTable[1][85] ) );
  LHQD1BWP \vrf/regTable_reg[1][86]  ( .E(n3588), .D(\vrf/N104 ), .Q(
        \vrf/regTable[1][86] ) );
  LHQD1BWP \vrf/regTable_reg[1][87]  ( .E(n3588), .D(\vrf/N105 ), .Q(
        \vrf/regTable[1][87] ) );
  LHQD1BWP \vrf/regTable_reg[1][88]  ( .E(n3588), .D(\vrf/N106 ), .Q(
        \vrf/regTable[1][88] ) );
  LHQD1BWP \vrf/regTable_reg[1][89]  ( .E(n3588), .D(\vrf/N107 ), .Q(
        \vrf/regTable[1][89] ) );
  LHQD1BWP \vrf/regTable_reg[1][90]  ( .E(n3588), .D(\vrf/N108 ), .Q(
        \vrf/regTable[1][90] ) );
  LHQD1BWP \vrf/regTable_reg[1][91]  ( .E(n3588), .D(\vrf/N109 ), .Q(
        \vrf/regTable[1][91] ) );
  LHQD1BWP \vrf/regTable_reg[1][92]  ( .E(n3588), .D(\vrf/N110 ), .Q(
        \vrf/regTable[1][92] ) );
  LHQD1BWP \vrf/regTable_reg[1][93]  ( .E(n3588), .D(\vrf/N111 ), .Q(
        \vrf/regTable[1][93] ) );
  LHQD1BWP \vrf/regTable_reg[1][94]  ( .E(n3588), .D(\vrf/N112 ), .Q(
        \vrf/regTable[1][94] ) );
  LHQD1BWP \vrf/regTable_reg[1][95]  ( .E(n3588), .D(\vrf/N113 ), .Q(
        \vrf/regTable[1][95] ) );
  LHQD1BWP \vrf/regTable_reg[1][96]  ( .E(n3588), .D(\vrf/N114 ), .Q(
        \vrf/regTable[1][96] ) );
  LHQD1BWP \vrf/regTable_reg[1][97]  ( .E(n3588), .D(\vrf/N115 ), .Q(
        \vrf/regTable[1][97] ) );
  LHQD1BWP \vrf/regTable_reg[1][98]  ( .E(n3588), .D(\vrf/N116 ), .Q(
        \vrf/regTable[1][98] ) );
  LHQD1BWP \vrf/regTable_reg[1][99]  ( .E(n3588), .D(\vrf/N118 ), .Q(
        \vrf/regTable[1][99] ) );
  LHQD1BWP \vrf/regTable_reg[1][100]  ( .E(n3588), .D(\vrf/N119 ), .Q(
        \vrf/regTable[1][100] ) );
  LHQD1BWP \vrf/regTable_reg[1][101]  ( .E(n3588), .D(\vrf/N120 ), .Q(
        \vrf/regTable[1][101] ) );
  LHQD1BWP \vrf/regTable_reg[1][102]  ( .E(n3588), .D(\vrf/N121 ), .Q(
        \vrf/regTable[1][102] ) );
  LHQD1BWP \vrf/regTable_reg[1][103]  ( .E(n3588), .D(\vrf/N122 ), .Q(
        \vrf/regTable[1][103] ) );
  LHQD1BWP \vrf/regTable_reg[1][104]  ( .E(n3588), .D(\vrf/N123 ), .Q(
        \vrf/regTable[1][104] ) );
  LHQD1BWP \vrf/regTable_reg[1][105]  ( .E(n3588), .D(\vrf/N124 ), .Q(
        \vrf/regTable[1][105] ) );
  LHQD1BWP \vrf/regTable_reg[1][106]  ( .E(n3588), .D(\vrf/N125 ), .Q(
        \vrf/regTable[1][106] ) );
  LHQD1BWP \vrf/regTable_reg[1][107]  ( .E(n3588), .D(\vrf/N126 ), .Q(
        \vrf/regTable[1][107] ) );
  LHQD1BWP \vrf/regTable_reg[1][108]  ( .E(n3588), .D(\vrf/N127 ), .Q(
        \vrf/regTable[1][108] ) );
  LHQD1BWP \vrf/regTable_reg[1][109]  ( .E(n3588), .D(\vrf/N128 ), .Q(
        \vrf/regTable[1][109] ) );
  LHQD1BWP \vrf/regTable_reg[1][110]  ( .E(n3588), .D(\vrf/N129 ), .Q(
        \vrf/regTable[1][110] ) );
  LHQD1BWP \vrf/regTable_reg[1][111]  ( .E(n3588), .D(\vrf/N130 ), .Q(
        \vrf/regTable[1][111] ) );
  LHQD1BWP \vrf/regTable_reg[1][112]  ( .E(n3588), .D(\vrf/N131 ), .Q(
        \vrf/regTable[1][112] ) );
  LHQD1BWP \vrf/regTable_reg[1][113]  ( .E(n3588), .D(\vrf/N132 ), .Q(
        \vrf/regTable[1][113] ) );
  LHQD1BWP \vrf/regTable_reg[1][114]  ( .E(n3588), .D(\vrf/N133 ), .Q(
        \vrf/regTable[1][114] ) );
  LHQD1BWP \vrf/regTable_reg[1][115]  ( .E(n3588), .D(\vrf/N134 ), .Q(
        \vrf/regTable[1][115] ) );
  LHQD1BWP \vrf/regTable_reg[1][116]  ( .E(n3588), .D(\vrf/N135 ), .Q(
        \vrf/regTable[1][116] ) );
  LHQD1BWP \vrf/regTable_reg[1][117]  ( .E(n3588), .D(\vrf/N136 ), .Q(
        \vrf/regTable[1][117] ) );
  LHQD1BWP \vrf/regTable_reg[1][118]  ( .E(n3588), .D(\vrf/N137 ), .Q(
        \vrf/regTable[1][118] ) );
  LHQD1BWP \vrf/regTable_reg[1][119]  ( .E(n3588), .D(\vrf/N138 ), .Q(
        \vrf/regTable[1][119] ) );
  LHQD1BWP \vrf/regTable_reg[1][120]  ( .E(n3588), .D(\vrf/N139 ), .Q(
        \vrf/regTable[1][120] ) );
  LHQD1BWP \vrf/regTable_reg[1][121]  ( .E(n3588), .D(\vrf/N140 ), .Q(
        \vrf/regTable[1][121] ) );
  LHQD1BWP \vrf/regTable_reg[1][122]  ( .E(n3588), .D(\vrf/N141 ), .Q(
        \vrf/regTable[1][122] ) );
  LHQD1BWP \vrf/regTable_reg[1][123]  ( .E(n3588), .D(\vrf/N142 ), .Q(
        \vrf/regTable[1][123] ) );
  LHQD1BWP \vrf/regTable_reg[1][124]  ( .E(n3588), .D(\vrf/N143 ), .Q(
        \vrf/regTable[1][124] ) );
  LHQD1BWP \vrf/regTable_reg[1][125]  ( .E(n3588), .D(\vrf/N144 ), .Q(
        \vrf/regTable[1][125] ) );
  LHQD1BWP \vrf/regTable_reg[1][126]  ( .E(n3588), .D(\vrf/N145 ), .Q(
        \vrf/regTable[1][126] ) );
  LHQD1BWP \vrf/regTable_reg[1][127]  ( .E(n3588), .D(\vrf/N146 ), .Q(
        \vrf/regTable[1][127] ) );
  LHQD1BWP \vrf/regTable_reg[1][128]  ( .E(n3588), .D(\vrf/N147 ), .Q(
        \vrf/regTable[1][128] ) );
  LHQD1BWP \vrf/regTable_reg[1][129]  ( .E(n3588), .D(\vrf/N148 ), .Q(
        \vrf/regTable[1][129] ) );
  LHQD1BWP \vrf/regTable_reg[1][130]  ( .E(n3588), .D(\vrf/N149 ), .Q(
        \vrf/regTable[1][130] ) );
  LHQD1BWP \vrf/regTable_reg[1][131]  ( .E(n3588), .D(\vrf/N150 ), .Q(
        \vrf/regTable[1][131] ) );
  LHQD1BWP \vrf/regTable_reg[1][132]  ( .E(n3588), .D(\vrf/N151 ), .Q(
        \vrf/regTable[1][132] ) );
  LHQD1BWP \vrf/regTable_reg[1][133]  ( .E(n3588), .D(\vrf/N152 ), .Q(
        \vrf/regTable[1][133] ) );
  LHQD1BWP \vrf/regTable_reg[1][134]  ( .E(n3588), .D(\vrf/N153 ), .Q(
        \vrf/regTable[1][134] ) );
  LHQD1BWP \vrf/regTable_reg[1][135]  ( .E(n3588), .D(\vrf/N154 ), .Q(
        \vrf/regTable[1][135] ) );
  LHQD1BWP \vrf/regTable_reg[1][136]  ( .E(n3588), .D(\vrf/N155 ), .Q(
        \vrf/regTable[1][136] ) );
  LHQD1BWP \vrf/regTable_reg[1][137]  ( .E(\vrf/N293 ), .D(\vrf/N156 ), .Q(
        \vrf/regTable[1][137] ) );
  LHQD1BWP \vrf/regTable_reg[1][138]  ( .E(n3588), .D(\vrf/N157 ), .Q(
        \vrf/regTable[1][138] ) );
  LHQD1BWP \vrf/regTable_reg[1][139]  ( .E(\vrf/N293 ), .D(\vrf/N158 ), .Q(
        \vrf/regTable[1][139] ) );
  LHQD1BWP \vrf/regTable_reg[1][140]  ( .E(n3588), .D(\vrf/N159 ), .Q(
        \vrf/regTable[1][140] ) );
  LHQD1BWP \vrf/regTable_reg[1][141]  ( .E(\vrf/N293 ), .D(\vrf/N160 ), .Q(
        \vrf/regTable[1][141] ) );
  LHQD1BWP \vrf/regTable_reg[1][142]  ( .E(n3588), .D(\vrf/N161 ), .Q(
        \vrf/regTable[1][142] ) );
  LHQD1BWP \vrf/regTable_reg[1][143]  ( .E(\vrf/N293 ), .D(\vrf/N162 ), .Q(
        \vrf/regTable[1][143] ) );
  LHQD1BWP \vrf/regTable_reg[1][144]  ( .E(n3588), .D(\vrf/N163 ), .Q(
        \vrf/regTable[1][144] ) );
  LHQD1BWP \vrf/regTable_reg[1][145]  ( .E(\vrf/N293 ), .D(\vrf/N164 ), .Q(
        \vrf/regTable[1][145] ) );
  LHQD1BWP \vrf/regTable_reg[1][146]  ( .E(n3588), .D(\vrf/N165 ), .Q(
        \vrf/regTable[1][146] ) );
  LHQD1BWP \vrf/regTable_reg[1][147]  ( .E(\vrf/N293 ), .D(\vrf/N166 ), .Q(
        \vrf/regTable[1][147] ) );
  LHQD1BWP \vrf/regTable_reg[1][148]  ( .E(n3588), .D(\vrf/N167 ), .Q(
        \vrf/regTable[1][148] ) );
  LHQD1BWP \vrf/regTable_reg[1][149]  ( .E(n3588), .D(\vrf/N168 ), .Q(
        \vrf/regTable[1][149] ) );
  LHQD1BWP \vrf/regTable_reg[1][150]  ( .E(n3588), .D(\vrf/N169 ), .Q(
        \vrf/regTable[1][150] ) );
  LHQD1BWP \vrf/regTable_reg[1][151]  ( .E(\vrf/N293 ), .D(\vrf/N170 ), .Q(
        \vrf/regTable[1][151] ) );
  LHQD1BWP \vrf/regTable_reg[1][152]  ( .E(n3588), .D(\vrf/N171 ), .Q(
        \vrf/regTable[1][152] ) );
  LHQD1BWP \vrf/regTable_reg[1][153]  ( .E(n3588), .D(\vrf/N172 ), .Q(
        \vrf/regTable[1][153] ) );
  LHQD1BWP \vrf/regTable_reg[1][154]  ( .E(n3588), .D(\vrf/N173 ), .Q(
        \vrf/regTable[1][154] ) );
  LHQD1BWP \vrf/regTable_reg[1][155]  ( .E(\vrf/N293 ), .D(\vrf/N174 ), .Q(
        \vrf/regTable[1][155] ) );
  LHQD1BWP \vrf/regTable_reg[1][156]  ( .E(n3588), .D(\vrf/N175 ), .Q(
        \vrf/regTable[1][156] ) );
  LHQD1BWP \vrf/regTable_reg[1][157]  ( .E(n3588), .D(\vrf/N176 ), .Q(
        \vrf/regTable[1][157] ) );
  LHQD1BWP \vrf/regTable_reg[1][158]  ( .E(n3588), .D(\vrf/N177 ), .Q(
        \vrf/regTable[1][158] ) );
  LHQD1BWP \vrf/regTable_reg[1][159]  ( .E(n3588), .D(\vrf/N178 ), .Q(
        \vrf/regTable[1][159] ) );
  LHQD1BWP \vrf/regTable_reg[1][160]  ( .E(\vrf/N293 ), .D(\vrf/N179 ), .Q(
        \vrf/regTable[1][160] ) );
  LHQD1BWP \vrf/regTable_reg[1][161]  ( .E(n3588), .D(\vrf/N180 ), .Q(
        \vrf/regTable[1][161] ) );
  LHQD1BWP \vrf/regTable_reg[1][162]  ( .E(n3588), .D(\vrf/N181 ), .Q(
        \vrf/regTable[1][162] ) );
  LHQD1BWP \vrf/regTable_reg[1][163]  ( .E(n3588), .D(\vrf/N182 ), .Q(
        \vrf/regTable[1][163] ) );
  LHQD1BWP \vrf/regTable_reg[1][164]  ( .E(\vrf/N293 ), .D(\vrf/N183 ), .Q(
        \vrf/regTable[1][164] ) );
  LHQD1BWP \vrf/regTable_reg[1][165]  ( .E(n3588), .D(\vrf/N184 ), .Q(
        \vrf/regTable[1][165] ) );
  LHQD1BWP \vrf/regTable_reg[1][166]  ( .E(n3588), .D(\vrf/N185 ), .Q(
        \vrf/regTable[1][166] ) );
  LHQD1BWP \vrf/regTable_reg[1][167]  ( .E(n3588), .D(\vrf/N186 ), .Q(
        \vrf/regTable[1][167] ) );
  LHQD1BWP \vrf/regTable_reg[1][168]  ( .E(\vrf/N293 ), .D(\vrf/N187 ), .Q(
        \vrf/regTable[1][168] ) );
  LHQD1BWP \vrf/regTable_reg[1][169]  ( .E(n3588), .D(\vrf/N188 ), .Q(
        \vrf/regTable[1][169] ) );
  LHQD1BWP \vrf/regTable_reg[1][170]  ( .E(n3588), .D(\vrf/N189 ), .Q(
        \vrf/regTable[1][170] ) );
  LHQD1BWP \vrf/regTable_reg[1][171]  ( .E(n3588), .D(\vrf/N190 ), .Q(
        \vrf/regTable[1][171] ) );
  LHQD1BWP \vrf/regTable_reg[1][172]  ( .E(n3588), .D(\vrf/N191 ), .Q(
        \vrf/regTable[1][172] ) );
  LHQD1BWP \vrf/regTable_reg[1][173]  ( .E(n3588), .D(\vrf/N192 ), .Q(
        \vrf/regTable[1][173] ) );
  LHQD1BWP \vrf/regTable_reg[1][174]  ( .E(\vrf/N293 ), .D(\vrf/N193 ), .Q(
        \vrf/regTable[1][174] ) );
  LHQD1BWP \vrf/regTable_reg[1][175]  ( .E(n3588), .D(\vrf/N194 ), .Q(
        \vrf/regTable[1][175] ) );
  LHQD1BWP \vrf/regTable_reg[1][176]  ( .E(n3588), .D(\vrf/N195 ), .Q(
        \vrf/regTable[1][176] ) );
  LHQD1BWP \vrf/regTable_reg[1][177]  ( .E(n3588), .D(\vrf/N196 ), .Q(
        \vrf/regTable[1][177] ) );
  LHQD1BWP \vrf/regTable_reg[1][178]  ( .E(n3588), .D(\vrf/N197 ), .Q(
        \vrf/regTable[1][178] ) );
  LHQD1BWP \vrf/regTable_reg[1][179]  ( .E(\vrf/N293 ), .D(\vrf/N198 ), .Q(
        \vrf/regTable[1][179] ) );
  LHQD1BWP \vrf/regTable_reg[1][180]  ( .E(n3588), .D(\vrf/N199 ), .Q(
        \vrf/regTable[1][180] ) );
  LHQD1BWP \vrf/regTable_reg[1][181]  ( .E(n3588), .D(\vrf/N200 ), .Q(
        \vrf/regTable[1][181] ) );
  LHQD1BWP \vrf/regTable_reg[1][182]  ( .E(n3588), .D(\vrf/N201 ), .Q(
        \vrf/regTable[1][182] ) );
  LHQD1BWP \vrf/regTable_reg[1][183]  ( .E(n3588), .D(\vrf/N202 ), .Q(
        \vrf/regTable[1][183] ) );
  LHQD1BWP \vrf/regTable_reg[1][184]  ( .E(n3588), .D(\vrf/N203 ), .Q(
        \vrf/regTable[1][184] ) );
  LHQD1BWP \vrf/regTable_reg[1][185]  ( .E(n3588), .D(\vrf/N204 ), .Q(
        \vrf/regTable[1][185] ) );
  LHQD1BWP \vrf/regTable_reg[1][186]  ( .E(n3588), .D(\vrf/N205 ), .Q(
        \vrf/regTable[1][186] ) );
  LHQD1BWP \vrf/regTable_reg[1][187]  ( .E(n3588), .D(\vrf/N206 ), .Q(
        \vrf/regTable[1][187] ) );
  LHQD1BWP \vrf/regTable_reg[1][188]  ( .E(n3588), .D(\vrf/N207 ), .Q(
        \vrf/regTable[1][188] ) );
  LHQD1BWP \vrf/regTable_reg[1][189]  ( .E(\vrf/N293 ), .D(\vrf/N208 ), .Q(
        \vrf/regTable[1][189] ) );
  LHQD1BWP \vrf/regTable_reg[1][190]  ( .E(n3588), .D(\vrf/N209 ), .Q(
        \vrf/regTable[1][190] ) );
  LHQD1BWP \vrf/regTable_reg[1][191]  ( .E(n3588), .D(\vrf/N210 ), .Q(
        \vrf/regTable[1][191] ) );
  LHQD1BWP \vrf/regTable_reg[1][192]  ( .E(n3588), .D(\vrf/N211 ), .Q(
        \vrf/regTable[1][192] ) );
  LHQD1BWP \vrf/regTable_reg[1][193]  ( .E(n3588), .D(\vrf/N212 ), .Q(
        \vrf/regTable[1][193] ) );
  LHQD1BWP \vrf/regTable_reg[1][194]  ( .E(\vrf/N293 ), .D(\vrf/N213 ), .Q(
        \vrf/regTable[1][194] ) );
  LHQD1BWP \vrf/regTable_reg[1][195]  ( .E(\vrf/N293 ), .D(\vrf/N214 ), .Q(
        \vrf/regTable[1][195] ) );
  LHQD1BWP \vrf/regTable_reg[1][196]  ( .E(n3588), .D(\vrf/N215 ), .Q(
        \vrf/regTable[1][196] ) );
  LHQD1BWP \vrf/regTable_reg[1][197]  ( .E(n3588), .D(\vrf/N216 ), .Q(
        \vrf/regTable[1][197] ) );
  LHQD1BWP \vrf/regTable_reg[1][198]  ( .E(n3588), .D(\vrf/N218 ), .Q(
        \vrf/regTable[1][198] ) );
  LHQD1BWP \vrf/regTable_reg[1][199]  ( .E(n3588), .D(\vrf/N219 ), .Q(
        \vrf/regTable[1][199] ) );
  LHQD1BWP \vrf/regTable_reg[1][200]  ( .E(n3588), .D(\vrf/N220 ), .Q(
        \vrf/regTable[1][200] ) );
  LHQD1BWP \vrf/regTable_reg[1][201]  ( .E(\vrf/N293 ), .D(\vrf/N221 ), .Q(
        \vrf/regTable[1][201] ) );
  LHQD1BWP \vrf/regTable_reg[1][202]  ( .E(n3588), .D(\vrf/N222 ), .Q(
        \vrf/regTable[1][202] ) );
  LHQD1BWP \vrf/regTable_reg[1][203]  ( .E(n3588), .D(\vrf/N223 ), .Q(
        \vrf/regTable[1][203] ) );
  LHQD1BWP \vrf/regTable_reg[1][204]  ( .E(\vrf/N293 ), .D(\vrf/N224 ), .Q(
        \vrf/regTable[1][204] ) );
  LHQD1BWP \vrf/regTable_reg[1][205]  ( .E(n3588), .D(\vrf/N225 ), .Q(
        \vrf/regTable[1][205] ) );
  LHQD1BWP \vrf/regTable_reg[1][206]  ( .E(\vrf/N293 ), .D(\vrf/N226 ), .Q(
        \vrf/regTable[1][206] ) );
  LHQD1BWP \vrf/regTable_reg[1][207]  ( .E(n3588), .D(\vrf/N227 ), .Q(
        \vrf/regTable[1][207] ) );
  LHQD1BWP \vrf/regTable_reg[1][208]  ( .E(n3588), .D(\vrf/N228 ), .Q(
        \vrf/regTable[1][208] ) );
  LHQD1BWP \vrf/regTable_reg[1][209]  ( .E(n3588), .D(\vrf/N229 ), .Q(
        \vrf/regTable[1][209] ) );
  LHQD1BWP \vrf/regTable_reg[1][210]  ( .E(n3588), .D(\vrf/N230 ), .Q(
        \vrf/regTable[1][210] ) );
  LHQD1BWP \vrf/regTable_reg[1][211]  ( .E(n3588), .D(\vrf/N231 ), .Q(
        \vrf/regTable[1][211] ) );
  LHQD1BWP \vrf/regTable_reg[1][212]  ( .E(n3588), .D(\vrf/N232 ), .Q(
        \vrf/regTable[1][212] ) );
  LHQD1BWP \vrf/regTable_reg[1][213]  ( .E(n3588), .D(\vrf/N233 ), .Q(
        \vrf/regTable[1][213] ) );
  LHQD1BWP \vrf/regTable_reg[1][214]  ( .E(n3588), .D(\vrf/N234 ), .Q(
        \vrf/regTable[1][214] ) );
  LHQD1BWP \vrf/regTable_reg[1][215]  ( .E(n3588), .D(\vrf/N235 ), .Q(
        \vrf/regTable[1][215] ) );
  LHQD1BWP \vrf/regTable_reg[1][216]  ( .E(n3588), .D(\vrf/N236 ), .Q(
        \vrf/regTable[1][216] ) );
  LHQD1BWP \vrf/regTable_reg[1][217]  ( .E(n3588), .D(\vrf/N237 ), .Q(
        \vrf/regTable[1][217] ) );
  LHQD1BWP \vrf/regTable_reg[1][218]  ( .E(n3588), .D(\vrf/N238 ), .Q(
        \vrf/regTable[1][218] ) );
  LHQD1BWP \vrf/regTable_reg[1][219]  ( .E(n3588), .D(\vrf/N239 ), .Q(
        \vrf/regTable[1][219] ) );
  LHQD1BWP \vrf/regTable_reg[1][220]  ( .E(n3588), .D(\vrf/N240 ), .Q(
        \vrf/regTable[1][220] ) );
  LHQD1BWP \vrf/regTable_reg[1][221]  ( .E(n3588), .D(\vrf/N241 ), .Q(
        \vrf/regTable[1][221] ) );
  LHQD1BWP \vrf/regTable_reg[1][222]  ( .E(n3588), .D(\vrf/N242 ), .Q(
        \vrf/regTable[1][222] ) );
  LHQD1BWP \vrf/regTable_reg[1][223]  ( .E(\vrf/N293 ), .D(\vrf/N243 ), .Q(
        \vrf/regTable[1][223] ) );
  LHQD1BWP \vrf/regTable_reg[1][224]  ( .E(n3588), .D(\vrf/N244 ), .Q(
        \vrf/regTable[1][224] ) );
  LHQD1BWP \vrf/regTable_reg[1][225]  ( .E(n3588), .D(\vrf/N245 ), .Q(
        \vrf/regTable[1][225] ) );
  LHQD1BWP \vrf/regTable_reg[1][226]  ( .E(n3588), .D(\vrf/N246 ), .Q(
        \vrf/regTable[1][226] ) );
  LHQD1BWP \vrf/regTable_reg[1][227]  ( .E(\vrf/N293 ), .D(\vrf/N247 ), .Q(
        \vrf/regTable[1][227] ) );
  LHQD1BWP \vrf/regTable_reg[1][228]  ( .E(n3588), .D(\vrf/N248 ), .Q(
        \vrf/regTable[1][228] ) );
  LHQD1BWP \vrf/regTable_reg[1][229]  ( .E(n3588), .D(\vrf/N249 ), .Q(
        \vrf/regTable[1][229] ) );
  LHQD1BWP \vrf/regTable_reg[1][230]  ( .E(n3588), .D(\vrf/N250 ), .Q(
        \vrf/regTable[1][230] ) );
  LHQD1BWP \vrf/regTable_reg[1][231]  ( .E(\vrf/N293 ), .D(\vrf/N251 ), .Q(
        \vrf/regTable[1][231] ) );
  LHQD1BWP \vrf/regTable_reg[1][232]  ( .E(n3588), .D(\vrf/N252 ), .Q(
        \vrf/regTable[1][232] ) );
  LHQD1BWP \vrf/regTable_reg[1][233]  ( .E(n3588), .D(\vrf/N253 ), .Q(
        \vrf/regTable[1][233] ) );
  LHQD1BWP \vrf/regTable_reg[1][234]  ( .E(n3588), .D(\vrf/N254 ), .Q(
        \vrf/regTable[1][234] ) );
  LHQD1BWP \vrf/regTable_reg[1][235]  ( .E(n3588), .D(\vrf/N255 ), .Q(
        \vrf/regTable[1][235] ) );
  LHQD1BWP \vrf/regTable_reg[1][236]  ( .E(n3588), .D(\vrf/N256 ), .Q(
        \vrf/regTable[1][236] ) );
  LHQD1BWP \vrf/regTable_reg[1][237]  ( .E(n3588), .D(\vrf/N257 ), .Q(
        \vrf/regTable[1][237] ) );
  LHQD1BWP \vrf/regTable_reg[1][238]  ( .E(n3588), .D(\vrf/N258 ), .Q(
        \vrf/regTable[1][238] ) );
  LHQD1BWP \vrf/regTable_reg[1][239]  ( .E(n3588), .D(\vrf/N259 ), .Q(
        \vrf/regTable[1][239] ) );
  LHQD1BWP \vrf/regTable_reg[1][240]  ( .E(n3588), .D(\vrf/N260 ), .Q(
        \vrf/regTable[1][240] ) );
  LHQD1BWP \vrf/regTable_reg[1][241]  ( .E(n3588), .D(\vrf/N261 ), .Q(
        \vrf/regTable[1][241] ) );
  LHQD1BWP \vrf/regTable_reg[1][242]  ( .E(n3588), .D(\vrf/N262 ), .Q(
        \vrf/regTable[1][242] ) );
  LHQD1BWP \vrf/regTable_reg[1][243]  ( .E(n3588), .D(\vrf/N263 ), .Q(
        \vrf/regTable[1][243] ) );
  LHQD1BWP \vrf/regTable_reg[1][244]  ( .E(n3588), .D(\vrf/N264 ), .Q(
        \vrf/regTable[1][244] ) );
  LHQD1BWP \vrf/regTable_reg[1][245]  ( .E(n3588), .D(\vrf/N265 ), .Q(
        \vrf/regTable[1][245] ) );
  LHQD1BWP \vrf/regTable_reg[1][246]  ( .E(n3588), .D(\vrf/N266 ), .Q(
        \vrf/regTable[1][246] ) );
  LHQD1BWP \vrf/regTable_reg[1][247]  ( .E(n3588), .D(\vrf/N267 ), .Q(
        \vrf/regTable[1][247] ) );
  LHQD1BWP \vrf/regTable_reg[1][248]  ( .E(n3588), .D(\vrf/N268 ), .Q(
        \vrf/regTable[1][248] ) );
  LHQD1BWP \vrf/regTable_reg[1][249]  ( .E(n3588), .D(\vrf/N269 ), .Q(
        \vrf/regTable[1][249] ) );
  LHQD1BWP \vrf/regTable_reg[1][250]  ( .E(n3588), .D(\vrf/N270 ), .Q(
        \vrf/regTable[1][250] ) );
  LHQD1BWP \vrf/regTable_reg[1][251]  ( .E(\vrf/N293 ), .D(\vrf/N271 ), .Q(
        \vrf/regTable[1][251] ) );
  LHQD1BWP \vrf/regTable_reg[1][252]  ( .E(n3588), .D(\vrf/N272 ), .Q(
        \vrf/regTable[1][252] ) );
  LHQD1BWP \vrf/regTable_reg[1][253]  ( .E(n3588), .D(\vrf/N273 ), .Q(
        \vrf/regTable[1][253] ) );
  LHQD1BWP \vrf/regTable_reg[1][254]  ( .E(n3588), .D(\vrf/N274 ), .Q(
        \vrf/regTable[1][254] ) );
  LHQD1BWP \vrf/regTable_reg[1][255]  ( .E(n3588), .D(\vrf/N275 ), .Q(
        \vrf/regTable[1][255] ) );
  LHQD1BWP \vrf/regTable_reg[0][0]  ( .E(n3590), .D(\vrf/N18 ), .Q(
        \vrf/regTable[0][0] ) );
  LHQD1BWP \vrf/regTable_reg[0][1]  ( .E(n3590), .D(\vrf/N19 ), .Q(
        \vrf/regTable[0][1] ) );
  LHQD1BWP \vrf/regTable_reg[0][2]  ( .E(n3590), .D(\vrf/N20 ), .Q(
        \vrf/regTable[0][2] ) );
  LHQD1BWP \vrf/regTable_reg[0][3]  ( .E(n3590), .D(\vrf/N21 ), .Q(
        \vrf/regTable[0][3] ) );
  LHQD1BWP \vrf/regTable_reg[0][4]  ( .E(n3590), .D(\vrf/N22 ), .Q(
        \vrf/regTable[0][4] ) );
  LHQD1BWP \vrf/regTable_reg[0][5]  ( .E(n3590), .D(\vrf/N23 ), .Q(
        \vrf/regTable[0][5] ) );
  LHQD1BWP \vrf/regTable_reg[0][6]  ( .E(n3590), .D(\vrf/N24 ), .Q(
        \vrf/regTable[0][6] ) );
  LHQD1BWP \vrf/regTable_reg[0][7]  ( .E(n3590), .D(\vrf/N25 ), .Q(
        \vrf/regTable[0][7] ) );
  LHQD1BWP \vrf/regTable_reg[0][8]  ( .E(n3590), .D(\vrf/N26 ), .Q(
        \vrf/regTable[0][8] ) );
  LHQD1BWP \vrf/regTable_reg[0][9]  ( .E(n3590), .D(\vrf/N27 ), .Q(
        \vrf/regTable[0][9] ) );
  LHQD1BWP \vrf/regTable_reg[0][10]  ( .E(n3590), .D(\vrf/N28 ), .Q(
        \vrf/regTable[0][10] ) );
  LHQD1BWP \vrf/regTable_reg[0][11]  ( .E(n3590), .D(\vrf/N29 ), .Q(
        \vrf/regTable[0][11] ) );
  LHQD1BWP \vrf/regTable_reg[0][12]  ( .E(n3590), .D(\vrf/N30 ), .Q(
        \vrf/regTable[0][12] ) );
  LHQD1BWP \vrf/regTable_reg[0][13]  ( .E(n3590), .D(\vrf/N31 ), .Q(
        \vrf/regTable[0][13] ) );
  LHQD1BWP \vrf/regTable_reg[0][14]  ( .E(n3590), .D(\vrf/N32 ), .Q(
        \vrf/regTable[0][14] ) );
  LHQD1BWP \vrf/regTable_reg[0][15]  ( .E(n3590), .D(\vrf/N33 ), .Q(
        \vrf/regTable[0][15] ) );
  LHQD1BWP \vrf/regTable_reg[0][16]  ( .E(n3590), .D(\vrf/N34 ), .Q(
        \vrf/regTable[0][16] ) );
  LHQD1BWP \vrf/regTable_reg[0][17]  ( .E(n3590), .D(\vrf/N35 ), .Q(
        \vrf/regTable[0][17] ) );
  LHQD1BWP \vrf/regTable_reg[0][18]  ( .E(n3590), .D(\vrf/N36 ), .Q(
        \vrf/regTable[0][18] ) );
  LHQD1BWP \vrf/regTable_reg[0][19]  ( .E(n3590), .D(\vrf/N37 ), .Q(
        \vrf/regTable[0][19] ) );
  LHQD1BWP \vrf/regTable_reg[0][20]  ( .E(n3590), .D(\vrf/N38 ), .Q(
        \vrf/regTable[0][20] ) );
  LHQD1BWP \vrf/regTable_reg[0][21]  ( .E(n3590), .D(\vrf/N39 ), .Q(
        \vrf/regTable[0][21] ) );
  LHQD1BWP \vrf/regTable_reg[0][22]  ( .E(n3590), .D(\vrf/N40 ), .Q(
        \vrf/regTable[0][22] ) );
  LHQD1BWP \vrf/regTable_reg[0][23]  ( .E(n3590), .D(\vrf/N41 ), .Q(
        \vrf/regTable[0][23] ) );
  LHQD1BWP \vrf/regTable_reg[0][24]  ( .E(n3590), .D(\vrf/N42 ), .Q(
        \vrf/regTable[0][24] ) );
  LHQD1BWP \vrf/regTable_reg[0][25]  ( .E(n3590), .D(\vrf/N43 ), .Q(
        \vrf/regTable[0][25] ) );
  LHQD1BWP \vrf/regTable_reg[0][26]  ( .E(n3590), .D(\vrf/N44 ), .Q(
        \vrf/regTable[0][26] ) );
  LHQD1BWP \vrf/regTable_reg[0][27]  ( .E(n3590), .D(\vrf/N45 ), .Q(
        \vrf/regTable[0][27] ) );
  LHQD1BWP \vrf/regTable_reg[0][28]  ( .E(n3590), .D(\vrf/N46 ), .Q(
        \vrf/regTable[0][28] ) );
  LHQD1BWP \vrf/regTable_reg[0][29]  ( .E(n3590), .D(\vrf/N47 ), .Q(
        \vrf/regTable[0][29] ) );
  LHQD1BWP \vrf/regTable_reg[0][30]  ( .E(n3590), .D(\vrf/N48 ), .Q(
        \vrf/regTable[0][30] ) );
  LHQD1BWP \vrf/regTable_reg[0][31]  ( .E(n3590), .D(\vrf/N49 ), .Q(
        \vrf/regTable[0][31] ) );
  LHQD1BWP \vrf/regTable_reg[0][32]  ( .E(n3590), .D(\vrf/N50 ), .Q(
        \vrf/regTable[0][32] ) );
  LHQD1BWP \vrf/regTable_reg[0][33]  ( .E(n3590), .D(\vrf/N51 ), .Q(
        \vrf/regTable[0][33] ) );
  LHQD1BWP \vrf/regTable_reg[0][34]  ( .E(n3590), .D(\vrf/N52 ), .Q(
        \vrf/regTable[0][34] ) );
  LHQD1BWP \vrf/regTable_reg[0][35]  ( .E(n3590), .D(\vrf/N53 ), .Q(
        \vrf/regTable[0][35] ) );
  LHQD1BWP \vrf/regTable_reg[0][36]  ( .E(n3590), .D(\vrf/N54 ), .Q(
        \vrf/regTable[0][36] ) );
  LHQD1BWP \vrf/regTable_reg[0][37]  ( .E(n3590), .D(\vrf/N55 ), .Q(
        \vrf/regTable[0][37] ) );
  LHQD1BWP \vrf/regTable_reg[0][38]  ( .E(n3590), .D(\vrf/N56 ), .Q(
        \vrf/regTable[0][38] ) );
  LHQD1BWP \vrf/regTable_reg[0][39]  ( .E(n3590), .D(\vrf/N57 ), .Q(
        \vrf/regTable[0][39] ) );
  LHQD1BWP \vrf/regTable_reg[0][40]  ( .E(n3590), .D(\vrf/N58 ), .Q(
        \vrf/regTable[0][40] ) );
  LHQD1BWP \vrf/regTable_reg[0][41]  ( .E(n3590), .D(\vrf/N59 ), .Q(
        \vrf/regTable[0][41] ) );
  LHQD1BWP \vrf/regTable_reg[0][42]  ( .E(n3590), .D(\vrf/N60 ), .Q(
        \vrf/regTable[0][42] ) );
  LHQD1BWP \vrf/regTable_reg[0][43]  ( .E(n3590), .D(\vrf/N61 ), .Q(
        \vrf/regTable[0][43] ) );
  LHQD1BWP \vrf/regTable_reg[0][44]  ( .E(n3590), .D(\vrf/N62 ), .Q(
        \vrf/regTable[0][44] ) );
  LHQD1BWP \vrf/regTable_reg[0][45]  ( .E(n3590), .D(\vrf/N63 ), .Q(
        \vrf/regTable[0][45] ) );
  LHQD1BWP \vrf/regTable_reg[0][46]  ( .E(n3590), .D(\vrf/N64 ), .Q(
        \vrf/regTable[0][46] ) );
  LHQD1BWP \vrf/regTable_reg[0][47]  ( .E(n3590), .D(\vrf/N65 ), .Q(
        \vrf/regTable[0][47] ) );
  LHQD1BWP \vrf/regTable_reg[0][48]  ( .E(n3590), .D(\vrf/N66 ), .Q(
        \vrf/regTable[0][48] ) );
  LHQD1BWP \vrf/regTable_reg[0][49]  ( .E(n3590), .D(\vrf/N67 ), .Q(
        \vrf/regTable[0][49] ) );
  LHQD1BWP \vrf/regTable_reg[0][50]  ( .E(n3590), .D(\vrf/N68 ), .Q(
        \vrf/regTable[0][50] ) );
  LHQD1BWP \vrf/regTable_reg[0][51]  ( .E(n3590), .D(\vrf/N69 ), .Q(
        \vrf/regTable[0][51] ) );
  LHQD1BWP \vrf/regTable_reg[0][52]  ( .E(n3590), .D(\vrf/N70 ), .Q(
        \vrf/regTable[0][52] ) );
  LHQD1BWP \vrf/regTable_reg[0][53]  ( .E(n3590), .D(\vrf/N71 ), .Q(
        \vrf/regTable[0][53] ) );
  LHQD1BWP \vrf/regTable_reg[0][54]  ( .E(n3590), .D(\vrf/N72 ), .Q(
        \vrf/regTable[0][54] ) );
  LHQD1BWP \vrf/regTable_reg[0][55]  ( .E(n3590), .D(\vrf/N73 ), .Q(
        \vrf/regTable[0][55] ) );
  LHQD1BWP \vrf/regTable_reg[0][56]  ( .E(n3590), .D(\vrf/N74 ), .Q(
        \vrf/regTable[0][56] ) );
  LHQD1BWP \vrf/regTable_reg[0][57]  ( .E(n3590), .D(\vrf/N75 ), .Q(
        \vrf/regTable[0][57] ) );
  LHQD1BWP \vrf/regTable_reg[0][58]  ( .E(n3590), .D(\vrf/N76 ), .Q(
        \vrf/regTable[0][58] ) );
  LHQD1BWP \vrf/regTable_reg[0][59]  ( .E(n3590), .D(\vrf/N77 ), .Q(
        \vrf/regTable[0][59] ) );
  LHQD1BWP \vrf/regTable_reg[0][60]  ( .E(n3590), .D(\vrf/N78 ), .Q(
        \vrf/regTable[0][60] ) );
  LHQD1BWP \vrf/regTable_reg[0][61]  ( .E(n3590), .D(\vrf/N79 ), .Q(
        \vrf/regTable[0][61] ) );
  LHQD1BWP \vrf/regTable_reg[0][62]  ( .E(n3590), .D(\vrf/N80 ), .Q(
        \vrf/regTable[0][62] ) );
  LHQD1BWP \vrf/regTable_reg[0][63]  ( .E(n3590), .D(\vrf/N81 ), .Q(
        \vrf/regTable[0][63] ) );
  LHQD1BWP \vrf/regTable_reg[0][64]  ( .E(n3590), .D(\vrf/N82 ), .Q(
        \vrf/regTable[0][64] ) );
  LHQD1BWP \vrf/regTable_reg[0][65]  ( .E(n3590), .D(\vrf/N83 ), .Q(
        \vrf/regTable[0][65] ) );
  LHQD1BWP \vrf/regTable_reg[0][66]  ( .E(n3590), .D(\vrf/N84 ), .Q(
        \vrf/regTable[0][66] ) );
  LHQD1BWP \vrf/regTable_reg[0][67]  ( .E(n3590), .D(\vrf/N85 ), .Q(
        \vrf/regTable[0][67] ) );
  LHQD1BWP \vrf/regTable_reg[0][68]  ( .E(n3590), .D(\vrf/N86 ), .Q(
        \vrf/regTable[0][68] ) );
  LHQD1BWP \vrf/regTable_reg[0][69]  ( .E(n3590), .D(\vrf/N87 ), .Q(
        \vrf/regTable[0][69] ) );
  LHQD1BWP \vrf/regTable_reg[0][70]  ( .E(n3590), .D(\vrf/N88 ), .Q(
        \vrf/regTable[0][70] ) );
  LHQD1BWP \vrf/regTable_reg[0][71]  ( .E(n3590), .D(\vrf/N89 ), .Q(
        \vrf/regTable[0][71] ) );
  LHQD1BWP \vrf/regTable_reg[0][72]  ( .E(n3590), .D(\vrf/N90 ), .Q(
        \vrf/regTable[0][72] ) );
  LHQD1BWP \vrf/regTable_reg[0][73]  ( .E(n3590), .D(\vrf/N91 ), .Q(
        \vrf/regTable[0][73] ) );
  LHQD1BWP \vrf/regTable_reg[0][74]  ( .E(n3590), .D(\vrf/N92 ), .Q(
        \vrf/regTable[0][74] ) );
  LHQD1BWP \vrf/regTable_reg[0][75]  ( .E(n3590), .D(\vrf/N93 ), .Q(
        \vrf/regTable[0][75] ) );
  LHQD1BWP \vrf/regTable_reg[0][76]  ( .E(n3590), .D(\vrf/N94 ), .Q(
        \vrf/regTable[0][76] ) );
  LHQD1BWP \vrf/regTable_reg[0][77]  ( .E(n3590), .D(\vrf/N95 ), .Q(
        \vrf/regTable[0][77] ) );
  LHQD1BWP \vrf/regTable_reg[0][78]  ( .E(n3590), .D(\vrf/N96 ), .Q(
        \vrf/regTable[0][78] ) );
  LHQD1BWP \vrf/regTable_reg[0][79]  ( .E(n3590), .D(\vrf/N97 ), .Q(
        \vrf/regTable[0][79] ) );
  LHQD1BWP \vrf/regTable_reg[0][80]  ( .E(n3590), .D(\vrf/N98 ), .Q(
        \vrf/regTable[0][80] ) );
  LHQD1BWP \vrf/regTable_reg[0][81]  ( .E(n3590), .D(\vrf/N99 ), .Q(
        \vrf/regTable[0][81] ) );
  LHQD1BWP \vrf/regTable_reg[0][82]  ( .E(n3590), .D(\vrf/N100 ), .Q(
        \vrf/regTable[0][82] ) );
  LHQD1BWP \vrf/regTable_reg[0][83]  ( .E(n3590), .D(\vrf/N101 ), .Q(
        \vrf/regTable[0][83] ) );
  LHQD1BWP \vrf/regTable_reg[0][84]  ( .E(n3590), .D(\vrf/N102 ), .Q(
        \vrf/regTable[0][84] ) );
  LHQD1BWP \vrf/regTable_reg[0][85]  ( .E(n3590), .D(\vrf/N103 ), .Q(
        \vrf/regTable[0][85] ) );
  LHQD1BWP \vrf/regTable_reg[0][86]  ( .E(n3590), .D(\vrf/N104 ), .Q(
        \vrf/regTable[0][86] ) );
  LHQD1BWP \vrf/regTable_reg[0][87]  ( .E(n3590), .D(\vrf/N105 ), .Q(
        \vrf/regTable[0][87] ) );
  LHQD1BWP \vrf/regTable_reg[0][88]  ( .E(n3590), .D(\vrf/N106 ), .Q(
        \vrf/regTable[0][88] ) );
  LHQD1BWP \vrf/regTable_reg[0][89]  ( .E(n3590), .D(\vrf/N107 ), .Q(
        \vrf/regTable[0][89] ) );
  LHQD1BWP \vrf/regTable_reg[0][90]  ( .E(n3590), .D(\vrf/N108 ), .Q(
        \vrf/regTable[0][90] ) );
  LHQD1BWP \vrf/regTable_reg[0][91]  ( .E(n3590), .D(\vrf/N109 ), .Q(
        \vrf/regTable[0][91] ) );
  LHQD1BWP \vrf/regTable_reg[0][92]  ( .E(n3590), .D(\vrf/N110 ), .Q(
        \vrf/regTable[0][92] ) );
  LHQD1BWP \vrf/regTable_reg[0][93]  ( .E(n3590), .D(\vrf/N111 ), .Q(
        \vrf/regTable[0][93] ) );
  LHQD1BWP \vrf/regTable_reg[0][94]  ( .E(n3590), .D(\vrf/N112 ), .Q(
        \vrf/regTable[0][94] ) );
  LHQD1BWP \vrf/regTable_reg[0][95]  ( .E(n3590), .D(\vrf/N113 ), .Q(
        \vrf/regTable[0][95] ) );
  LHQD1BWP \vrf/regTable_reg[0][96]  ( .E(n3590), .D(\vrf/N114 ), .Q(
        \vrf/regTable[0][96] ) );
  LHQD1BWP \vrf/regTable_reg[0][97]  ( .E(n3590), .D(\vrf/N115 ), .Q(
        \vrf/regTable[0][97] ) );
  LHQD1BWP \vrf/regTable_reg[0][98]  ( .E(n3590), .D(\vrf/N116 ), .Q(
        \vrf/regTable[0][98] ) );
  LHQD1BWP \vrf/regTable_reg[0][99]  ( .E(n3590), .D(\vrf/N118 ), .Q(
        \vrf/regTable[0][99] ) );
  LHQD1BWP \vrf/regTable_reg[0][100]  ( .E(n3590), .D(\vrf/N119 ), .Q(
        \vrf/regTable[0][100] ) );
  LHQD1BWP \vrf/regTable_reg[0][101]  ( .E(n3590), .D(\vrf/N120 ), .Q(
        \vrf/regTable[0][101] ) );
  LHQD1BWP \vrf/regTable_reg[0][102]  ( .E(n3590), .D(\vrf/N121 ), .Q(
        \vrf/regTable[0][102] ) );
  LHQD1BWP \vrf/regTable_reg[0][103]  ( .E(n3590), .D(\vrf/N122 ), .Q(
        \vrf/regTable[0][103] ) );
  LHQD1BWP \vrf/regTable_reg[0][104]  ( .E(n3590), .D(\vrf/N123 ), .Q(
        \vrf/regTable[0][104] ) );
  LHQD1BWP \vrf/regTable_reg[0][105]  ( .E(n3590), .D(\vrf/N124 ), .Q(
        \vrf/regTable[0][105] ) );
  LHQD1BWP \vrf/regTable_reg[0][106]  ( .E(n3590), .D(\vrf/N125 ), .Q(
        \vrf/regTable[0][106] ) );
  LHQD1BWP \vrf/regTable_reg[0][107]  ( .E(n3590), .D(\vrf/N126 ), .Q(
        \vrf/regTable[0][107] ) );
  LHQD1BWP \vrf/regTable_reg[0][108]  ( .E(n3590), .D(\vrf/N127 ), .Q(
        \vrf/regTable[0][108] ) );
  LHQD1BWP \vrf/regTable_reg[0][109]  ( .E(n3590), .D(\vrf/N128 ), .Q(
        \vrf/regTable[0][109] ) );
  LHQD1BWP \vrf/regTable_reg[0][110]  ( .E(n3590), .D(\vrf/N129 ), .Q(
        \vrf/regTable[0][110] ) );
  LHQD1BWP \vrf/regTable_reg[0][111]  ( .E(n3590), .D(\vrf/N130 ), .Q(
        \vrf/regTable[0][111] ) );
  LHQD1BWP \vrf/regTable_reg[0][112]  ( .E(n3590), .D(\vrf/N131 ), .Q(
        \vrf/regTable[0][112] ) );
  LHQD1BWP \vrf/regTable_reg[0][113]  ( .E(n3590), .D(\vrf/N132 ), .Q(
        \vrf/regTable[0][113] ) );
  LHQD1BWP \vrf/regTable_reg[0][114]  ( .E(n3590), .D(\vrf/N133 ), .Q(
        \vrf/regTable[0][114] ) );
  LHQD1BWP \vrf/regTable_reg[0][115]  ( .E(n3590), .D(\vrf/N134 ), .Q(
        \vrf/regTable[0][115] ) );
  LHQD1BWP \vrf/regTable_reg[0][116]  ( .E(n3590), .D(\vrf/N135 ), .Q(
        \vrf/regTable[0][116] ) );
  LHQD1BWP \vrf/regTable_reg[0][117]  ( .E(n3590), .D(\vrf/N136 ), .Q(
        \vrf/regTable[0][117] ) );
  LHQD1BWP \vrf/regTable_reg[0][118]  ( .E(n3590), .D(\vrf/N137 ), .Q(
        \vrf/regTable[0][118] ) );
  LHQD1BWP \vrf/regTable_reg[0][119]  ( .E(n3590), .D(\vrf/N138 ), .Q(
        \vrf/regTable[0][119] ) );
  LHQD1BWP \vrf/regTable_reg[0][120]  ( .E(n3590), .D(\vrf/N139 ), .Q(
        \vrf/regTable[0][120] ) );
  LHQD1BWP \vrf/regTable_reg[0][121]  ( .E(n3590), .D(\vrf/N140 ), .Q(
        \vrf/regTable[0][121] ) );
  LHQD1BWP \vrf/regTable_reg[0][122]  ( .E(n3590), .D(\vrf/N141 ), .Q(
        \vrf/regTable[0][122] ) );
  LHQD1BWP \vrf/regTable_reg[0][123]  ( .E(n3590), .D(\vrf/N142 ), .Q(
        \vrf/regTable[0][123] ) );
  LHQD1BWP \vrf/regTable_reg[0][124]  ( .E(n3590), .D(\vrf/N143 ), .Q(
        \vrf/regTable[0][124] ) );
  LHQD1BWP \vrf/regTable_reg[0][125]  ( .E(n3590), .D(\vrf/N144 ), .Q(
        \vrf/regTable[0][125] ) );
  LHQD1BWP \vrf/regTable_reg[0][126]  ( .E(n3590), .D(\vrf/N145 ), .Q(
        \vrf/regTable[0][126] ) );
  LHQD1BWP \vrf/regTable_reg[0][127]  ( .E(n3590), .D(\vrf/N146 ), .Q(
        \vrf/regTable[0][127] ) );
  LHQD1BWP \vrf/regTable_reg[0][128]  ( .E(n3590), .D(\vrf/N147 ), .Q(
        \vrf/regTable[0][128] ) );
  LHQD1BWP \vrf/regTable_reg[0][129]  ( .E(n3590), .D(\vrf/N148 ), .Q(
        \vrf/regTable[0][129] ) );
  LHQD1BWP \vrf/regTable_reg[0][130]  ( .E(n3590), .D(\vrf/N149 ), .Q(
        \vrf/regTable[0][130] ) );
  LHQD1BWP \vrf/regTable_reg[0][131]  ( .E(n3590), .D(\vrf/N150 ), .Q(
        \vrf/regTable[0][131] ) );
  LHQD1BWP \vrf/regTable_reg[0][132]  ( .E(n3590), .D(\vrf/N151 ), .Q(
        \vrf/regTable[0][132] ) );
  LHQD1BWP \vrf/regTable_reg[0][133]  ( .E(n3590), .D(\vrf/N152 ), .Q(
        \vrf/regTable[0][133] ) );
  LHQD1BWP \vrf/regTable_reg[0][134]  ( .E(n3590), .D(\vrf/N153 ), .Q(
        \vrf/regTable[0][134] ) );
  LHQD1BWP \vrf/regTable_reg[0][135]  ( .E(n3590), .D(\vrf/N154 ), .Q(
        \vrf/regTable[0][135] ) );
  LHQD1BWP \vrf/regTable_reg[0][136]  ( .E(n3590), .D(\vrf/N155 ), .Q(
        \vrf/regTable[0][136] ) );
  LHQD1BWP \vrf/regTable_reg[0][137]  ( .E(\vrf/N296 ), .D(\vrf/N156 ), .Q(
        \vrf/regTable[0][137] ) );
  LHQD1BWP \vrf/regTable_reg[0][138]  ( .E(n3590), .D(\vrf/N157 ), .Q(
        \vrf/regTable[0][138] ) );
  LHQD1BWP \vrf/regTable_reg[0][139]  ( .E(\vrf/N296 ), .D(\vrf/N158 ), .Q(
        \vrf/regTable[0][139] ) );
  LHQD1BWP \vrf/regTable_reg[0][140]  ( .E(n3590), .D(\vrf/N159 ), .Q(
        \vrf/regTable[0][140] ) );
  LHQD1BWP \vrf/regTable_reg[0][141]  ( .E(\vrf/N296 ), .D(\vrf/N160 ), .Q(
        \vrf/regTable[0][141] ) );
  LHQD1BWP \vrf/regTable_reg[0][142]  ( .E(n3590), .D(\vrf/N161 ), .Q(
        \vrf/regTable[0][142] ) );
  LHQD1BWP \vrf/regTable_reg[0][143]  ( .E(\vrf/N296 ), .D(\vrf/N162 ), .Q(
        \vrf/regTable[0][143] ) );
  LHQD1BWP \vrf/regTable_reg[0][144]  ( .E(n3590), .D(\vrf/N163 ), .Q(
        \vrf/regTable[0][144] ) );
  LHQD1BWP \vrf/regTable_reg[0][145]  ( .E(\vrf/N296 ), .D(\vrf/N164 ), .Q(
        \vrf/regTable[0][145] ) );
  LHQD1BWP \vrf/regTable_reg[0][146]  ( .E(n3590), .D(\vrf/N165 ), .Q(
        \vrf/regTable[0][146] ) );
  LHQD1BWP \vrf/regTable_reg[0][147]  ( .E(\vrf/N296 ), .D(\vrf/N166 ), .Q(
        \vrf/regTable[0][147] ) );
  LHQD1BWP \vrf/regTable_reg[0][148]  ( .E(n3590), .D(\vrf/N167 ), .Q(
        \vrf/regTable[0][148] ) );
  LHQD1BWP \vrf/regTable_reg[0][149]  ( .E(n3590), .D(\vrf/N168 ), .Q(
        \vrf/regTable[0][149] ) );
  LHQD1BWP \vrf/regTable_reg[0][150]  ( .E(n3590), .D(\vrf/N169 ), .Q(
        \vrf/regTable[0][150] ) );
  LHQD1BWP \vrf/regTable_reg[0][151]  ( .E(\vrf/N296 ), .D(\vrf/N170 ), .Q(
        \vrf/regTable[0][151] ) );
  LHQD1BWP \vrf/regTable_reg[0][152]  ( .E(n3590), .D(\vrf/N171 ), .Q(
        \vrf/regTable[0][152] ) );
  LHQD1BWP \vrf/regTable_reg[0][153]  ( .E(n3590), .D(\vrf/N172 ), .Q(
        \vrf/regTable[0][153] ) );
  LHQD1BWP \vrf/regTable_reg[0][154]  ( .E(n3590), .D(\vrf/N173 ), .Q(
        \vrf/regTable[0][154] ) );
  LHQD1BWP \vrf/regTable_reg[0][155]  ( .E(\vrf/N296 ), .D(\vrf/N174 ), .Q(
        \vrf/regTable[0][155] ) );
  LHQD1BWP \vrf/regTable_reg[0][156]  ( .E(n3590), .D(\vrf/N175 ), .Q(
        \vrf/regTable[0][156] ) );
  LHQD1BWP \vrf/regTable_reg[0][157]  ( .E(n3590), .D(\vrf/N176 ), .Q(
        \vrf/regTable[0][157] ) );
  LHQD1BWP \vrf/regTable_reg[0][158]  ( .E(n3590), .D(\vrf/N177 ), .Q(
        \vrf/regTable[0][158] ) );
  LHQD1BWP \vrf/regTable_reg[0][159]  ( .E(n3590), .D(\vrf/N178 ), .Q(
        \vrf/regTable[0][159] ) );
  LHQD1BWP \vrf/regTable_reg[0][160]  ( .E(\vrf/N296 ), .D(\vrf/N179 ), .Q(
        \vrf/regTable[0][160] ) );
  LHQD1BWP \vrf/regTable_reg[0][161]  ( .E(n3590), .D(\vrf/N180 ), .Q(
        \vrf/regTable[0][161] ) );
  LHQD1BWP \vrf/regTable_reg[0][162]  ( .E(n3590), .D(\vrf/N181 ), .Q(
        \vrf/regTable[0][162] ) );
  LHQD1BWP \vrf/regTable_reg[0][163]  ( .E(n3590), .D(\vrf/N182 ), .Q(
        \vrf/regTable[0][163] ) );
  LHQD1BWP \vrf/regTable_reg[0][164]  ( .E(\vrf/N296 ), .D(\vrf/N183 ), .Q(
        \vrf/regTable[0][164] ) );
  LHQD1BWP \vrf/regTable_reg[0][165]  ( .E(n3590), .D(\vrf/N184 ), .Q(
        \vrf/regTable[0][165] ) );
  LHQD1BWP \vrf/regTable_reg[0][166]  ( .E(n3590), .D(\vrf/N185 ), .Q(
        \vrf/regTable[0][166] ) );
  LHQD1BWP \vrf/regTable_reg[0][167]  ( .E(n3590), .D(\vrf/N186 ), .Q(
        \vrf/regTable[0][167] ) );
  LHQD1BWP \vrf/regTable_reg[0][168]  ( .E(\vrf/N296 ), .D(\vrf/N187 ), .Q(
        \vrf/regTable[0][168] ) );
  LHQD1BWP \vrf/regTable_reg[0][169]  ( .E(n3590), .D(\vrf/N188 ), .Q(
        \vrf/regTable[0][169] ) );
  LHQD1BWP \vrf/regTable_reg[0][170]  ( .E(n3590), .D(\vrf/N189 ), .Q(
        \vrf/regTable[0][170] ) );
  LHQD1BWP \vrf/regTable_reg[0][171]  ( .E(n3590), .D(\vrf/N190 ), .Q(
        \vrf/regTable[0][171] ) );
  LHQD1BWP \vrf/regTable_reg[0][172]  ( .E(n3590), .D(\vrf/N191 ), .Q(
        \vrf/regTable[0][172] ) );
  LHQD1BWP \vrf/regTable_reg[0][173]  ( .E(n3590), .D(\vrf/N192 ), .Q(
        \vrf/regTable[0][173] ) );
  LHQD1BWP \vrf/regTable_reg[0][174]  ( .E(\vrf/N296 ), .D(\vrf/N193 ), .Q(
        \vrf/regTable[0][174] ) );
  LHQD1BWP \vrf/regTable_reg[0][175]  ( .E(n3590), .D(\vrf/N194 ), .Q(
        \vrf/regTable[0][175] ) );
  LHQD1BWP \vrf/regTable_reg[0][176]  ( .E(n3590), .D(\vrf/N195 ), .Q(
        \vrf/regTable[0][176] ) );
  LHQD1BWP \vrf/regTable_reg[0][177]  ( .E(n3590), .D(\vrf/N196 ), .Q(
        \vrf/regTable[0][177] ) );
  LHQD1BWP \vrf/regTable_reg[0][178]  ( .E(n3590), .D(\vrf/N197 ), .Q(
        \vrf/regTable[0][178] ) );
  LHQD1BWP \vrf/regTable_reg[0][179]  ( .E(\vrf/N296 ), .D(\vrf/N198 ), .Q(
        \vrf/regTable[0][179] ) );
  LHQD1BWP \vrf/regTable_reg[0][180]  ( .E(n3590), .D(\vrf/N199 ), .Q(
        \vrf/regTable[0][180] ) );
  LHQD1BWP \vrf/regTable_reg[0][181]  ( .E(n3590), .D(\vrf/N200 ), .Q(
        \vrf/regTable[0][181] ) );
  LHQD1BWP \vrf/regTable_reg[0][182]  ( .E(n3590), .D(\vrf/N201 ), .Q(
        \vrf/regTable[0][182] ) );
  LHQD1BWP \vrf/regTable_reg[0][183]  ( .E(n3590), .D(\vrf/N202 ), .Q(
        \vrf/regTable[0][183] ) );
  LHQD1BWP \vrf/regTable_reg[0][184]  ( .E(n3590), .D(\vrf/N203 ), .Q(
        \vrf/regTable[0][184] ) );
  LHQD1BWP \vrf/regTable_reg[0][185]  ( .E(n3590), .D(\vrf/N204 ), .Q(
        \vrf/regTable[0][185] ) );
  LHQD1BWP \vrf/regTable_reg[0][186]  ( .E(n3590), .D(\vrf/N205 ), .Q(
        \vrf/regTable[0][186] ) );
  LHQD1BWP \vrf/regTable_reg[0][187]  ( .E(n3590), .D(\vrf/N206 ), .Q(
        \vrf/regTable[0][187] ) );
  LHQD1BWP \vrf/regTable_reg[0][188]  ( .E(n3590), .D(\vrf/N207 ), .Q(
        \vrf/regTable[0][188] ) );
  LHQD1BWP \vrf/regTable_reg[0][189]  ( .E(\vrf/N296 ), .D(\vrf/N208 ), .Q(
        \vrf/regTable[0][189] ) );
  LHQD1BWP \vrf/regTable_reg[0][190]  ( .E(n3590), .D(\vrf/N209 ), .Q(
        \vrf/regTable[0][190] ) );
  LHQD1BWP \vrf/regTable_reg[0][191]  ( .E(n3590), .D(\vrf/N210 ), .Q(
        \vrf/regTable[0][191] ) );
  LHQD1BWP \vrf/regTable_reg[0][192]  ( .E(n3590), .D(\vrf/N211 ), .Q(
        \vrf/regTable[0][192] ) );
  LHQD1BWP \vrf/regTable_reg[0][193]  ( .E(n3590), .D(\vrf/N212 ), .Q(
        \vrf/regTable[0][193] ) );
  LHQD1BWP \vrf/regTable_reg[0][194]  ( .E(\vrf/N296 ), .D(\vrf/N213 ), .Q(
        \vrf/regTable[0][194] ) );
  LHQD1BWP \vrf/regTable_reg[0][195]  ( .E(\vrf/N296 ), .D(\vrf/N214 ), .Q(
        \vrf/regTable[0][195] ) );
  LHQD1BWP \vrf/regTable_reg[0][196]  ( .E(n3590), .D(\vrf/N215 ), .Q(
        \vrf/regTable[0][196] ) );
  LHQD1BWP \vrf/regTable_reg[0][197]  ( .E(n3590), .D(\vrf/N216 ), .Q(
        \vrf/regTable[0][197] ) );
  LHQD1BWP \vrf/regTable_reg[0][198]  ( .E(n3590), .D(\vrf/N218 ), .Q(
        \vrf/regTable[0][198] ) );
  LHQD1BWP \vrf/regTable_reg[0][199]  ( .E(n3590), .D(\vrf/N219 ), .Q(
        \vrf/regTable[0][199] ) );
  LHQD1BWP \vrf/regTable_reg[0][200]  ( .E(n3590), .D(\vrf/N220 ), .Q(
        \vrf/regTable[0][200] ) );
  LHQD1BWP \vrf/regTable_reg[0][201]  ( .E(\vrf/N296 ), .D(\vrf/N221 ), .Q(
        \vrf/regTable[0][201] ) );
  LHQD1BWP \vrf/regTable_reg[0][202]  ( .E(n3590), .D(\vrf/N222 ), .Q(
        \vrf/regTable[0][202] ) );
  LHQD1BWP \vrf/regTable_reg[0][203]  ( .E(n3590), .D(\vrf/N223 ), .Q(
        \vrf/regTable[0][203] ) );
  LHQD1BWP \vrf/regTable_reg[0][204]  ( .E(\vrf/N296 ), .D(\vrf/N224 ), .Q(
        \vrf/regTable[0][204] ) );
  LHQD1BWP \vrf/regTable_reg[0][205]  ( .E(n3590), .D(\vrf/N225 ), .Q(
        \vrf/regTable[0][205] ) );
  LHQD1BWP \vrf/regTable_reg[0][206]  ( .E(\vrf/N296 ), .D(\vrf/N226 ), .Q(
        \vrf/regTable[0][206] ) );
  LHQD1BWP \vrf/regTable_reg[0][207]  ( .E(n3590), .D(\vrf/N227 ), .Q(
        \vrf/regTable[0][207] ) );
  LHQD1BWP \vrf/regTable_reg[0][208]  ( .E(n3590), .D(\vrf/N228 ), .Q(
        \vrf/regTable[0][208] ) );
  LHQD1BWP \vrf/regTable_reg[0][209]  ( .E(n3590), .D(\vrf/N229 ), .Q(
        \vrf/regTable[0][209] ) );
  LHQD1BWP \vrf/regTable_reg[0][210]  ( .E(n3590), .D(\vrf/N230 ), .Q(
        \vrf/regTable[0][210] ) );
  LHQD1BWP \vrf/regTable_reg[0][211]  ( .E(n3590), .D(\vrf/N231 ), .Q(
        \vrf/regTable[0][211] ) );
  LHQD1BWP \vrf/regTable_reg[0][212]  ( .E(n3590), .D(\vrf/N232 ), .Q(
        \vrf/regTable[0][212] ) );
  LHQD1BWP \vrf/regTable_reg[0][213]  ( .E(n3590), .D(\vrf/N233 ), .Q(
        \vrf/regTable[0][213] ) );
  LHQD1BWP \vrf/regTable_reg[0][214]  ( .E(n3590), .D(\vrf/N234 ), .Q(
        \vrf/regTable[0][214] ) );
  LHQD1BWP \vrf/regTable_reg[0][215]  ( .E(n3590), .D(\vrf/N235 ), .Q(
        \vrf/regTable[0][215] ) );
  LHQD1BWP \vrf/regTable_reg[0][216]  ( .E(n3590), .D(\vrf/N236 ), .Q(
        \vrf/regTable[0][216] ) );
  LHQD1BWP \vrf/regTable_reg[0][217]  ( .E(n3590), .D(\vrf/N237 ), .Q(
        \vrf/regTable[0][217] ) );
  LHQD1BWP \vrf/regTable_reg[0][218]  ( .E(n3590), .D(\vrf/N238 ), .Q(
        \vrf/regTable[0][218] ) );
  LHQD1BWP \vrf/regTable_reg[0][219]  ( .E(n3590), .D(\vrf/N239 ), .Q(
        \vrf/regTable[0][219] ) );
  LHQD1BWP \vrf/regTable_reg[0][220]  ( .E(n3590), .D(\vrf/N240 ), .Q(
        \vrf/regTable[0][220] ) );
  LHQD1BWP \vrf/regTable_reg[0][221]  ( .E(n3590), .D(\vrf/N241 ), .Q(
        \vrf/regTable[0][221] ) );
  LHQD1BWP \vrf/regTable_reg[0][222]  ( .E(n3590), .D(\vrf/N242 ), .Q(
        \vrf/regTable[0][222] ) );
  LHQD1BWP \vrf/regTable_reg[0][223]  ( .E(\vrf/N296 ), .D(\vrf/N243 ), .Q(
        \vrf/regTable[0][223] ) );
  LHQD1BWP \vrf/regTable_reg[0][224]  ( .E(n3590), .D(\vrf/N244 ), .Q(
        \vrf/regTable[0][224] ) );
  LHQD1BWP \vrf/regTable_reg[0][225]  ( .E(n3590), .D(\vrf/N245 ), .Q(
        \vrf/regTable[0][225] ) );
  LHQD1BWP \vrf/regTable_reg[0][226]  ( .E(n3590), .D(\vrf/N246 ), .Q(
        \vrf/regTable[0][226] ) );
  LHQD1BWP \vrf/regTable_reg[0][227]  ( .E(\vrf/N296 ), .D(\vrf/N247 ), .Q(
        \vrf/regTable[0][227] ) );
  LHQD1BWP \vrf/regTable_reg[0][228]  ( .E(n3590), .D(\vrf/N248 ), .Q(
        \vrf/regTable[0][228] ) );
  LHQD1BWP \vrf/regTable_reg[0][229]  ( .E(n3590), .D(\vrf/N249 ), .Q(
        \vrf/regTable[0][229] ) );
  LHQD1BWP \vrf/regTable_reg[0][230]  ( .E(n3590), .D(\vrf/N250 ), .Q(
        \vrf/regTable[0][230] ) );
  LHQD1BWP \vrf/regTable_reg[0][231]  ( .E(\vrf/N296 ), .D(\vrf/N251 ), .Q(
        \vrf/regTable[0][231] ) );
  LHQD1BWP \vrf/regTable_reg[0][232]  ( .E(n3590), .D(\vrf/N252 ), .Q(
        \vrf/regTable[0][232] ) );
  LHQD1BWP \vrf/regTable_reg[0][233]  ( .E(n3590), .D(\vrf/N253 ), .Q(
        \vrf/regTable[0][233] ) );
  LHQD1BWP \vrf/regTable_reg[0][234]  ( .E(n3590), .D(\vrf/N254 ), .Q(
        \vrf/regTable[0][234] ) );
  LHQD1BWP \vrf/regTable_reg[0][235]  ( .E(n3590), .D(\vrf/N255 ), .Q(
        \vrf/regTable[0][235] ) );
  LHQD1BWP \vrf/regTable_reg[0][236]  ( .E(n3590), .D(\vrf/N256 ), .Q(
        \vrf/regTable[0][236] ) );
  LHQD1BWP \vrf/regTable_reg[0][237]  ( .E(n3590), .D(\vrf/N257 ), .Q(
        \vrf/regTable[0][237] ) );
  LHQD1BWP \vrf/regTable_reg[0][238]  ( .E(n3590), .D(\vrf/N258 ), .Q(
        \vrf/regTable[0][238] ) );
  LHQD1BWP \vrf/regTable_reg[0][239]  ( .E(n3590), .D(\vrf/N259 ), .Q(
        \vrf/regTable[0][239] ) );
  LHQD1BWP \vrf/regTable_reg[0][240]  ( .E(n3590), .D(\vrf/N260 ), .Q(
        \vrf/regTable[0][240] ) );
  LHQD1BWP \vrf/regTable_reg[0][241]  ( .E(n3590), .D(\vrf/N261 ), .Q(
        \vrf/regTable[0][241] ) );
  LHQD1BWP \vrf/regTable_reg[0][242]  ( .E(n3590), .D(\vrf/N262 ), .Q(
        \vrf/regTable[0][242] ) );
  LHQD1BWP \vrf/regTable_reg[0][243]  ( .E(n3590), .D(\vrf/N263 ), .Q(
        \vrf/regTable[0][243] ) );
  LHQD1BWP \vrf/regTable_reg[0][244]  ( .E(n3590), .D(\vrf/N264 ), .Q(
        \vrf/regTable[0][244] ) );
  LHQD1BWP \vrf/regTable_reg[0][245]  ( .E(n3590), .D(\vrf/N265 ), .Q(
        \vrf/regTable[0][245] ) );
  LHQD1BWP \vrf/regTable_reg[0][246]  ( .E(n3590), .D(\vrf/N266 ), .Q(
        \vrf/regTable[0][246] ) );
  LHQD1BWP \vrf/regTable_reg[0][247]  ( .E(n3590), .D(\vrf/N267 ), .Q(
        \vrf/regTable[0][247] ) );
  LHQD1BWP \vrf/regTable_reg[0][248]  ( .E(n3590), .D(\vrf/N268 ), .Q(
        \vrf/regTable[0][248] ) );
  LHQD1BWP \vrf/regTable_reg[0][249]  ( .E(n3590), .D(\vrf/N269 ), .Q(
        \vrf/regTable[0][249] ) );
  LHQD1BWP \vrf/regTable_reg[0][250]  ( .E(n3590), .D(\vrf/N270 ), .Q(
        \vrf/regTable[0][250] ) );
  LHQD1BWP \vrf/regTable_reg[0][251]  ( .E(\vrf/N296 ), .D(\vrf/N271 ), .Q(
        \vrf/regTable[0][251] ) );
  LHQD1BWP \vrf/regTable_reg[0][252]  ( .E(n3590), .D(\vrf/N272 ), .Q(
        \vrf/regTable[0][252] ) );
  LHQD1BWP \vrf/regTable_reg[0][253]  ( .E(n3590), .D(\vrf/N273 ), .Q(
        \vrf/regTable[0][253] ) );
  LHQD1BWP \vrf/regTable_reg[0][254]  ( .E(n3590), .D(\vrf/N274 ), .Q(
        \vrf/regTable[0][254] ) );
  LHQD1BWP \vrf/regTable_reg[0][255]  ( .E(n3590), .D(\vrf/N275 ), .Q(
        \vrf/regTable[0][255] ) );
  LHQD1BWP \srf/regTable_reg[7][0]  ( .E(\srf/N36 ), .D(\srf/N37 ), .Q(
        \srf/regTable[7][0] ) );
  LHQD1BWP \srf/regTable_reg[7][1]  ( .E(\srf/N36 ), .D(\srf/N38 ), .Q(
        \srf/regTable[7][1] ) );
  LHQD1BWP \srf/regTable_reg[7][2]  ( .E(\srf/N36 ), .D(\srf/N39 ), .Q(
        \srf/regTable[7][2] ) );
  LHQD1BWP \srf/regTable_reg[7][3]  ( .E(\srf/N36 ), .D(\srf/N40 ), .Q(
        \srf/regTable[7][3] ) );
  LHQD1BWP \srf/regTable_reg[7][4]  ( .E(\srf/N36 ), .D(\srf/N41 ), .Q(
        \srf/regTable[7][4] ) );
  LHQD1BWP \srf/regTable_reg[7][5]  ( .E(\srf/N36 ), .D(\srf/N42 ), .Q(
        \srf/regTable[7][5] ) );
  LHQD1BWP \srf/regTable_reg[7][6]  ( .E(\srf/N36 ), .D(\srf/N43 ), .Q(
        \srf/regTable[7][6] ) );
  LHQD1BWP \srf/regTable_reg[7][7]  ( .E(\srf/N36 ), .D(\srf/N44 ), .Q(
        \srf/regTable[7][7] ) );
  LHQD1BWP \srf/regTable_reg[7][8]  ( .E(\srf/N36 ), .D(\srf/N45 ), .Q(
        \srf/regTable[7][8] ) );
  LHQD1BWP \srf/regTable_reg[7][9]  ( .E(\srf/N36 ), .D(\srf/N46 ), .Q(
        \srf/regTable[7][9] ) );
  LHQD1BWP \srf/regTable_reg[7][10]  ( .E(\srf/N36 ), .D(\srf/N47 ), .Q(
        \srf/regTable[7][10] ) );
  LHQD1BWP \srf/regTable_reg[7][11]  ( .E(\srf/N36 ), .D(\srf/N48 ), .Q(
        \srf/regTable[7][11] ) );
  LHQD1BWP \srf/regTable_reg[7][12]  ( .E(\srf/N36 ), .D(\srf/N49 ), .Q(
        \srf/regTable[7][12] ) );
  LHQD1BWP \srf/regTable_reg[7][13]  ( .E(\srf/N36 ), .D(\srf/N50 ), .Q(
        \srf/regTable[7][13] ) );
  LHQD1BWP \srf/regTable_reg[7][14]  ( .E(\srf/N36 ), .D(\srf/N51 ), .Q(
        \srf/regTable[7][14] ) );
  LHQD1BWP \srf/regTable_reg[7][15]  ( .E(\srf/N36 ), .D(\srf/N52 ), .Q(
        \srf/regTable[7][15] ) );
  LHQD1BWP \srf/regTable_reg[6][0]  ( .E(\srf/N53 ), .D(\srf/N37 ), .Q(
        \srf/regTable[6][0] ) );
  LHQD1BWP \srf/regTable_reg[6][1]  ( .E(\srf/N53 ), .D(\srf/N38 ), .Q(
        \srf/regTable[6][1] ) );
  LHQD1BWP \srf/regTable_reg[6][2]  ( .E(\srf/N53 ), .D(\srf/N39 ), .Q(
        \srf/regTable[6][2] ) );
  LHQD1BWP \srf/regTable_reg[6][3]  ( .E(\srf/N53 ), .D(\srf/N40 ), .Q(
        \srf/regTable[6][3] ) );
  LHQD1BWP \srf/regTable_reg[6][4]  ( .E(\srf/N53 ), .D(\srf/N41 ), .Q(
        \srf/regTable[6][4] ) );
  LHQD1BWP \srf/regTable_reg[6][5]  ( .E(\srf/N53 ), .D(\srf/N42 ), .Q(
        \srf/regTable[6][5] ) );
  LHQD1BWP \srf/regTable_reg[6][6]  ( .E(\srf/N53 ), .D(\srf/N43 ), .Q(
        \srf/regTable[6][6] ) );
  LHQD1BWP \srf/regTable_reg[6][7]  ( .E(\srf/N53 ), .D(\srf/N44 ), .Q(
        \srf/regTable[6][7] ) );
  LHQD1BWP \srf/regTable_reg[6][8]  ( .E(\srf/N53 ), .D(\srf/N45 ), .Q(
        \srf/regTable[6][8] ) );
  LHQD1BWP \srf/regTable_reg[6][9]  ( .E(\srf/N53 ), .D(\srf/N46 ), .Q(
        \srf/regTable[6][9] ) );
  LHQD1BWP \srf/regTable_reg[6][10]  ( .E(\srf/N53 ), .D(\srf/N47 ), .Q(
        \srf/regTable[6][10] ) );
  LHQD1BWP \srf/regTable_reg[6][11]  ( .E(\srf/N53 ), .D(\srf/N48 ), .Q(
        \srf/regTable[6][11] ) );
  LHQD1BWP \srf/regTable_reg[6][12]  ( .E(\srf/N53 ), .D(\srf/N49 ), .Q(
        \srf/regTable[6][12] ) );
  LHQD1BWP \srf/regTable_reg[6][13]  ( .E(\srf/N53 ), .D(\srf/N50 ), .Q(
        \srf/regTable[6][13] ) );
  LHQD1BWP \srf/regTable_reg[6][14]  ( .E(\srf/N53 ), .D(\srf/N51 ), .Q(
        \srf/regTable[6][14] ) );
  LHQD1BWP \srf/regTable_reg[6][15]  ( .E(\srf/N53 ), .D(\srf/N52 ), .Q(
        \srf/regTable[6][15] ) );
  LHQD1BWP \srf/regTable_reg[5][0]  ( .E(\srf/N54 ), .D(\srf/N37 ), .Q(
        \srf/regTable[5][0] ) );
  LHQD1BWP \srf/regTable_reg[5][1]  ( .E(\srf/N54 ), .D(\srf/N38 ), .Q(
        \srf/regTable[5][1] ) );
  LHQD1BWP \srf/regTable_reg[5][2]  ( .E(\srf/N54 ), .D(\srf/N39 ), .Q(
        \srf/regTable[5][2] ) );
  LHQD1BWP \srf/regTable_reg[5][3]  ( .E(\srf/N54 ), .D(\srf/N40 ), .Q(
        \srf/regTable[5][3] ) );
  LHQD1BWP \srf/regTable_reg[5][4]  ( .E(\srf/N54 ), .D(\srf/N41 ), .Q(
        \srf/regTable[5][4] ) );
  LHQD1BWP \srf/regTable_reg[5][5]  ( .E(\srf/N54 ), .D(\srf/N42 ), .Q(
        \srf/regTable[5][5] ) );
  LHQD1BWP \srf/regTable_reg[5][6]  ( .E(\srf/N54 ), .D(\srf/N43 ), .Q(
        \srf/regTable[5][6] ) );
  LHQD1BWP \srf/regTable_reg[5][7]  ( .E(\srf/N54 ), .D(\srf/N44 ), .Q(
        \srf/regTable[5][7] ) );
  LHQD1BWP \srf/regTable_reg[5][8]  ( .E(\srf/N54 ), .D(\srf/N45 ), .Q(
        \srf/regTable[5][8] ) );
  LHQD1BWP \srf/regTable_reg[5][9]  ( .E(\srf/N54 ), .D(\srf/N46 ), .Q(
        \srf/regTable[5][9] ) );
  LHQD1BWP \srf/regTable_reg[5][10]  ( .E(\srf/N54 ), .D(\srf/N47 ), .Q(
        \srf/regTable[5][10] ) );
  LHQD1BWP \srf/regTable_reg[5][11]  ( .E(\srf/N54 ), .D(\srf/N48 ), .Q(
        \srf/regTable[5][11] ) );
  LHQD1BWP \srf/regTable_reg[5][12]  ( .E(\srf/N54 ), .D(\srf/N49 ), .Q(
        \srf/regTable[5][12] ) );
  LHQD1BWP \srf/regTable_reg[5][13]  ( .E(\srf/N54 ), .D(\srf/N50 ), .Q(
        \srf/regTable[5][13] ) );
  LHQD1BWP \srf/regTable_reg[5][14]  ( .E(\srf/N54 ), .D(\srf/N51 ), .Q(
        \srf/regTable[5][14] ) );
  LHQD1BWP \srf/regTable_reg[5][15]  ( .E(\srf/N54 ), .D(\srf/N52 ), .Q(
        \srf/regTable[5][15] ) );
  LHQD1BWP \srf/regTable_reg[4][0]  ( .E(\srf/N55 ), .D(\srf/N37 ), .Q(
        \srf/regTable[4][0] ) );
  LHQD1BWP \srf/regTable_reg[4][1]  ( .E(\srf/N55 ), .D(\srf/N38 ), .Q(
        \srf/regTable[4][1] ) );
  LHQD1BWP \srf/regTable_reg[4][2]  ( .E(\srf/N55 ), .D(\srf/N39 ), .Q(
        \srf/regTable[4][2] ) );
  LHQD1BWP \srf/regTable_reg[4][3]  ( .E(\srf/N55 ), .D(\srf/N40 ), .Q(
        \srf/regTable[4][3] ) );
  LHQD1BWP \srf/regTable_reg[4][4]  ( .E(\srf/N55 ), .D(\srf/N41 ), .Q(
        \srf/regTable[4][4] ) );
  LHQD1BWP \srf/regTable_reg[4][5]  ( .E(\srf/N55 ), .D(\srf/N42 ), .Q(
        \srf/regTable[4][5] ) );
  LHQD1BWP \srf/regTable_reg[4][6]  ( .E(\srf/N55 ), .D(\srf/N43 ), .Q(
        \srf/regTable[4][6] ) );
  LHQD1BWP \srf/regTable_reg[4][7]  ( .E(\srf/N55 ), .D(\srf/N44 ), .Q(
        \srf/regTable[4][7] ) );
  LHQD1BWP \srf/regTable_reg[4][8]  ( .E(\srf/N55 ), .D(\srf/N45 ), .Q(
        \srf/regTable[4][8] ) );
  LHQD1BWP \srf/regTable_reg[4][9]  ( .E(\srf/N55 ), .D(\srf/N46 ), .Q(
        \srf/regTable[4][9] ) );
  LHQD1BWP \srf/regTable_reg[4][10]  ( .E(\srf/N55 ), .D(\srf/N47 ), .Q(
        \srf/regTable[4][10] ) );
  LHQD1BWP \srf/regTable_reg[4][11]  ( .E(\srf/N55 ), .D(\srf/N48 ), .Q(
        \srf/regTable[4][11] ) );
  LHQD1BWP \srf/regTable_reg[4][12]  ( .E(\srf/N55 ), .D(\srf/N49 ), .Q(
        \srf/regTable[4][12] ) );
  LHQD1BWP \srf/regTable_reg[4][13]  ( .E(\srf/N55 ), .D(\srf/N50 ), .Q(
        \srf/regTable[4][13] ) );
  LHQD1BWP \srf/regTable_reg[4][14]  ( .E(\srf/N55 ), .D(\srf/N51 ), .Q(
        \srf/regTable[4][14] ) );
  LHQD1BWP \srf/regTable_reg[4][15]  ( .E(\srf/N55 ), .D(\srf/N52 ), .Q(
        \srf/regTable[4][15] ) );
  LHQD1BWP \srf/regTable_reg[3][0]  ( .E(\srf/N56 ), .D(\srf/N37 ), .Q(
        \srf/regTable[3][0] ) );
  LHQD1BWP \srf/regTable_reg[3][1]  ( .E(\srf/N56 ), .D(\srf/N38 ), .Q(
        \srf/regTable[3][1] ) );
  LHQD1BWP \srf/regTable_reg[3][2]  ( .E(\srf/N56 ), .D(\srf/N39 ), .Q(
        \srf/regTable[3][2] ) );
  LHQD1BWP \srf/regTable_reg[3][3]  ( .E(\srf/N56 ), .D(\srf/N40 ), .Q(
        \srf/regTable[3][3] ) );
  LHQD1BWP \srf/regTable_reg[3][4]  ( .E(\srf/N56 ), .D(\srf/N41 ), .Q(
        \srf/regTable[3][4] ) );
  LHQD1BWP \srf/regTable_reg[3][5]  ( .E(\srf/N56 ), .D(\srf/N42 ), .Q(
        \srf/regTable[3][5] ) );
  LHQD1BWP \srf/regTable_reg[3][6]  ( .E(\srf/N56 ), .D(\srf/N43 ), .Q(
        \srf/regTable[3][6] ) );
  LHQD1BWP \srf/regTable_reg[3][7]  ( .E(\srf/N56 ), .D(\srf/N44 ), .Q(
        \srf/regTable[3][7] ) );
  LHQD1BWP \srf/regTable_reg[3][8]  ( .E(\srf/N56 ), .D(\srf/N45 ), .Q(
        \srf/regTable[3][8] ) );
  LHQD1BWP \srf/regTable_reg[3][9]  ( .E(\srf/N56 ), .D(\srf/N46 ), .Q(
        \srf/regTable[3][9] ) );
  LHQD1BWP \srf/regTable_reg[3][10]  ( .E(\srf/N56 ), .D(\srf/N47 ), .Q(
        \srf/regTable[3][10] ) );
  LHQD1BWP \srf/regTable_reg[3][11]  ( .E(\srf/N56 ), .D(\srf/N48 ), .Q(
        \srf/regTable[3][11] ) );
  LHQD1BWP \srf/regTable_reg[3][12]  ( .E(\srf/N56 ), .D(\srf/N49 ), .Q(
        \srf/regTable[3][12] ) );
  LHQD1BWP \srf/regTable_reg[3][13]  ( .E(\srf/N56 ), .D(\srf/N50 ), .Q(
        \srf/regTable[3][13] ) );
  LHQD1BWP \srf/regTable_reg[3][14]  ( .E(\srf/N56 ), .D(\srf/N51 ), .Q(
        \srf/regTable[3][14] ) );
  LHQD1BWP \srf/regTable_reg[3][15]  ( .E(\srf/N56 ), .D(\srf/N52 ), .Q(
        \srf/regTable[3][15] ) );
  LHQD1BWP \srf/regTable_reg[2][0]  ( .E(\srf/N57 ), .D(\srf/N37 ), .Q(
        \srf/regTable[2][0] ) );
  LHQD1BWP \srf/regTable_reg[2][1]  ( .E(\srf/N57 ), .D(\srf/N38 ), .Q(
        \srf/regTable[2][1] ) );
  LHQD1BWP \srf/regTable_reg[2][2]  ( .E(\srf/N57 ), .D(\srf/N39 ), .Q(
        \srf/regTable[2][2] ) );
  LHQD1BWP \srf/regTable_reg[2][3]  ( .E(\srf/N57 ), .D(\srf/N40 ), .Q(
        \srf/regTable[2][3] ) );
  LHQD1BWP \srf/regTable_reg[2][4]  ( .E(\srf/N57 ), .D(\srf/N41 ), .Q(
        \srf/regTable[2][4] ) );
  LHQD1BWP \srf/regTable_reg[2][5]  ( .E(\srf/N57 ), .D(\srf/N42 ), .Q(
        \srf/regTable[2][5] ) );
  LHQD1BWP \srf/regTable_reg[2][6]  ( .E(\srf/N57 ), .D(\srf/N43 ), .Q(
        \srf/regTable[2][6] ) );
  LHQD1BWP \srf/regTable_reg[2][7]  ( .E(\srf/N57 ), .D(\srf/N44 ), .Q(
        \srf/regTable[2][7] ) );
  LHQD1BWP \srf/regTable_reg[2][8]  ( .E(\srf/N57 ), .D(\srf/N45 ), .Q(
        \srf/regTable[2][8] ) );
  LHQD1BWP \srf/regTable_reg[2][9]  ( .E(\srf/N57 ), .D(\srf/N46 ), .Q(
        \srf/regTable[2][9] ) );
  LHQD1BWP \srf/regTable_reg[2][10]  ( .E(\srf/N57 ), .D(\srf/N47 ), .Q(
        \srf/regTable[2][10] ) );
  LHQD1BWP \srf/regTable_reg[2][11]  ( .E(\srf/N57 ), .D(\srf/N48 ), .Q(
        \srf/regTable[2][11] ) );
  LHQD1BWP \srf/regTable_reg[2][12]  ( .E(\srf/N57 ), .D(\srf/N49 ), .Q(
        \srf/regTable[2][12] ) );
  LHQD1BWP \srf/regTable_reg[2][13]  ( .E(\srf/N57 ), .D(\srf/N50 ), .Q(
        \srf/regTable[2][13] ) );
  LHQD1BWP \srf/regTable_reg[2][14]  ( .E(\srf/N57 ), .D(\srf/N51 ), .Q(
        \srf/regTable[2][14] ) );
  LHQD1BWP \srf/regTable_reg[2][15]  ( .E(\srf/N57 ), .D(\srf/N52 ), .Q(
        \srf/regTable[2][15] ) );
  LHQD1BWP \srf/regTable_reg[1][0]  ( .E(\srf/N58 ), .D(\srf/N37 ), .Q(
        \srf/regTable[1][0] ) );
  LHQD1BWP \srf/regTable_reg[1][1]  ( .E(\srf/N58 ), .D(\srf/N38 ), .Q(
        \srf/regTable[1][1] ) );
  LHQD1BWP \srf/regTable_reg[1][2]  ( .E(\srf/N58 ), .D(\srf/N39 ), .Q(
        \srf/regTable[1][2] ) );
  LHQD1BWP \srf/regTable_reg[1][3]  ( .E(\srf/N58 ), .D(\srf/N40 ), .Q(
        \srf/regTable[1][3] ) );
  LHQD1BWP \srf/regTable_reg[1][4]  ( .E(\srf/N58 ), .D(\srf/N41 ), .Q(
        \srf/regTable[1][4] ) );
  LHQD1BWP \srf/regTable_reg[1][5]  ( .E(\srf/N58 ), .D(\srf/N42 ), .Q(
        \srf/regTable[1][5] ) );
  LHQD1BWP \srf/regTable_reg[1][6]  ( .E(\srf/N58 ), .D(\srf/N43 ), .Q(
        \srf/regTable[1][6] ) );
  LHQD1BWP \srf/regTable_reg[1][7]  ( .E(\srf/N58 ), .D(\srf/N44 ), .Q(
        \srf/regTable[1][7] ) );
  LHQD1BWP \srf/regTable_reg[1][8]  ( .E(\srf/N58 ), .D(\srf/N45 ), .Q(
        \srf/regTable[1][8] ) );
  LHQD1BWP \srf/regTable_reg[1][9]  ( .E(\srf/N58 ), .D(\srf/N46 ), .Q(
        \srf/regTable[1][9] ) );
  LHQD1BWP \srf/regTable_reg[1][10]  ( .E(\srf/N58 ), .D(\srf/N47 ), .Q(
        \srf/regTable[1][10] ) );
  LHQD1BWP \srf/regTable_reg[1][11]  ( .E(\srf/N58 ), .D(\srf/N48 ), .Q(
        \srf/regTable[1][11] ) );
  LHQD1BWP \srf/regTable_reg[1][12]  ( .E(\srf/N58 ), .D(\srf/N49 ), .Q(
        \srf/regTable[1][12] ) );
  LHQD1BWP \srf/regTable_reg[1][13]  ( .E(\srf/N58 ), .D(\srf/N50 ), .Q(
        \srf/regTable[1][13] ) );
  LHQD1BWP \srf/regTable_reg[1][14]  ( .E(\srf/N58 ), .D(\srf/N51 ), .Q(
        \srf/regTable[1][14] ) );
  LHQD1BWP \srf/regTable_reg[1][15]  ( .E(\srf/N58 ), .D(\srf/N52 ), .Q(
        \srf/regTable[1][15] ) );
  LHQD1BWP \srf/regTable_reg[0][0]  ( .E(\srf/N59 ), .D(\srf/N37 ), .Q(
        \srf/regTable[0][0] ) );
  LHQD1BWP \srf/regTable_reg[0][1]  ( .E(\srf/N59 ), .D(\srf/N38 ), .Q(
        \srf/regTable[0][1] ) );
  LHQD1BWP \srf/regTable_reg[0][2]  ( .E(\srf/N59 ), .D(\srf/N39 ), .Q(
        \srf/regTable[0][2] ) );
  LHQD1BWP \srf/regTable_reg[0][3]  ( .E(\srf/N59 ), .D(\srf/N40 ), .Q(
        \srf/regTable[0][3] ) );
  LHQD1BWP \srf/regTable_reg[0][4]  ( .E(\srf/N59 ), .D(\srf/N41 ), .Q(
        \srf/regTable[0][4] ) );
  LHQD1BWP \srf/regTable_reg[0][5]  ( .E(\srf/N59 ), .D(\srf/N42 ), .Q(
        \srf/regTable[0][5] ) );
  LHQD1BWP \srf/regTable_reg[0][6]  ( .E(\srf/N59 ), .D(\srf/N43 ), .Q(
        \srf/regTable[0][6] ) );
  LHQD1BWP \srf/regTable_reg[0][7]  ( .E(\srf/N59 ), .D(\srf/N44 ), .Q(
        \srf/regTable[0][7] ) );
  LHQD1BWP \srf/regTable_reg[0][8]  ( .E(\srf/N59 ), .D(\srf/N45 ), .Q(
        \srf/regTable[0][8] ) );
  LHQD1BWP \srf/regTable_reg[0][9]  ( .E(\srf/N59 ), .D(\srf/N46 ), .Q(
        \srf/regTable[0][9] ) );
  LHQD1BWP \srf/regTable_reg[0][10]  ( .E(\srf/N59 ), .D(\srf/N47 ), .Q(
        \srf/regTable[0][10] ) );
  LHQD1BWP \srf/regTable_reg[0][11]  ( .E(\srf/N59 ), .D(\srf/N48 ), .Q(
        \srf/regTable[0][11] ) );
  LHQD1BWP \srf/regTable_reg[0][12]  ( .E(\srf/N59 ), .D(\srf/N49 ), .Q(
        \srf/regTable[0][12] ) );
  LHQD1BWP \srf/regTable_reg[0][13]  ( .E(\srf/N59 ), .D(\srf/N50 ), .Q(
        \srf/regTable[0][13] ) );
  LHQD1BWP \srf/regTable_reg[0][14]  ( .E(\srf/N59 ), .D(\srf/N51 ), .Q(
        \srf/regTable[0][14] ) );
  LHQD1BWP \srf/regTable_reg[0][15]  ( .E(\srf/N59 ), .D(\srf/N52 ), .Q(
        \srf/regTable[0][15] ) );
  CMPE42D1BWP \mult_x_153/U55  ( .A(\mult_x_153/n181 ), .B(\mult_x_153/n148 ), 
        .C(\mult_x_153/n159 ), .CIX(\mult_x_153/n105 ), .D(\mult_x_153/n170 ), 
        .CO(\mult_x_153/n101 ), .COX(\mult_x_153/n100 ), .S(\mult_x_153/n102 )
         );
  CMPE42D1BWP \mult_x_153/U53  ( .A(\mult_x_153/n158 ), .B(\mult_x_153/n180 ), 
        .C(\mult_x_153/n169 ), .CIX(\mult_x_153/n100 ), .D(\mult_x_153/n99 ), 
        .CO(\mult_x_153/n96 ), .COX(\mult_x_153/n95 ), .S(\mult_x_153/n97 ) );
  CMPE42D1BWP \mult_x_153/U51  ( .A(\mult_x_153/n168 ), .B(\mult_x_153/n179 ), 
        .C(\mult_x_153/n98 ), .CIX(\mult_x_153/n94 ), .D(\mult_x_153/n95 ), 
        .CO(\mult_x_153/n91 ), .COX(\mult_x_153/n90 ), .S(\mult_x_153/n92 ) );
  CMPE42D1BWP \mult_x_153/U48  ( .A(\mult_x_153/n89 ), .B(\mult_x_153/n178 ), 
        .C(\mult_x_153/n93 ), .CIX(\mult_x_153/n90 ), .D(\mult_x_153/n87 ), 
        .CO(\mult_x_153/n84 ), .COX(\mult_x_153/n83 ), .S(\mult_x_153/n85 ) );
  CMPE42D1BWP \mult_x_153/U47  ( .A(\mult_x_153/n144 ), .B(\mult_x_153/n122 ), 
        .C(\mult_x_153/n177 ), .CIX(\mult_x_153/n88 ), .D(\mult_x_153/n133 ), 
        .CO(\mult_x_153/n81 ), .COX(\mult_x_153/n80 ), .S(\mult_x_153/n82 ) );
  CMPE42D1BWP \mult_x_153/U46  ( .A(\mult_x_153/n155 ), .B(\mult_x_153/n166 ), 
        .C(\mult_x_153/n86 ), .CIX(\mult_x_153/n82 ), .D(\mult_x_153/n83 ), 
        .CO(\mult_x_153/n78 ), .COX(\mult_x_153/n77 ), .S(\mult_x_153/n79 ) );
  CMPE42D1BWP \mult_x_153/U45  ( .A(\mult_x_153/n143 ), .B(\mult_x_153/n121 ), 
        .C(\mult_x_153/n176 ), .CIX(\mult_x_153/n154 ), .D(\mult_x_153/n132 ), 
        .CO(\mult_x_153/n75 ), .COX(\mult_x_153/n74 ), .S(\mult_x_153/n76 ) );
  CMPE42D1BWP \mult_x_153/U44  ( .A(\mult_x_153/n80 ), .B(\mult_x_153/n165 ), 
        .C(\mult_x_153/n77 ), .CIX(\mult_x_153/n81 ), .D(\mult_x_153/n76 ), 
        .CO(\mult_x_153/n72 ), .COX(\mult_x_153/n71 ), .S(\mult_x_153/n73 ) );
  CMPE42D1BWP \mult_x_153/U42  ( .A(\mult_x_153/n142 ), .B(\mult_x_153/n70 ), 
        .C(\mult_x_153/n131 ), .CIX(\mult_x_153/n74 ), .D(n6070), .CO(
        \mult_x_153/n68 ), .COX(\mult_x_153/n67 ), .S(\mult_x_153/n69 ) );
  CMPE42D1BWP \mult_x_153/U41  ( .A(\mult_x_153/n153 ), .B(\mult_x_153/n164 ), 
        .C(\mult_x_153/n69 ), .CIX(\mult_x_153/n71 ), .D(\mult_x_153/n75 ), 
        .CO(\mult_x_153/n65 ), .COX(\mult_x_153/n64 ), .S(\mult_x_153/n66 ) );
  CMPE42D1BWP \mult_x_153/U39  ( .A(\mult_x_153/n70 ), .B(\mult_x_153/n120 ), 
        .C(\mult_x_153/n163 ), .CIX(\mult_x_153/n130 ), .D(\mult_x_153/n152 ), 
        .CO(\mult_x_153/n60 ), .COX(\mult_x_153/n59 ), .S(\mult_x_153/n61 ) );
  CMPE42D1BWP \mult_x_153/U38  ( .A(\mult_x_153/n67 ), .B(\mult_x_153/n141 ), 
        .C(\mult_x_153/n61 ), .CIX(\mult_x_153/n64 ), .D(\mult_x_153/n68 ), 
        .CO(\mult_x_153/n57 ), .COX(\mult_x_153/n56 ), .S(\mult_x_153/n58 ) );
  CMPE42D1BWP \mult_x_153/U37  ( .A(\mult_x_153/n119 ), .B(n6071), .C(
        \mult_x_153/n151 ), .CIX(\mult_x_153/n59 ), .D(\mult_x_153/n162 ), 
        .CO(\mult_x_153/n54 ), .COX(\mult_x_153/n53 ), .S(\mult_x_153/n55 ) );
  CMPE42D1BWP \mult_x_153/U36  ( .A(\mult_x_153/n129 ), .B(\mult_x_153/n140 ), 
        .C(\mult_x_153/n55 ), .CIX(\mult_x_153/n56 ), .D(\mult_x_153/n60 ), 
        .CO(\mult_x_153/n51 ), .COX(\mult_x_153/n50 ), .S(\mult_x_153/n52 ) );
  CMPE42D1BWP \mult_x_153/U33  ( .A(\mult_x_153/n53 ), .B(\mult_x_153/n150 ), 
        .C(\mult_x_153/n47 ), .CIX(\mult_x_153/n50 ), .D(\mult_x_153/n54 ), 
        .CO(\mult_x_153/n44 ), .COX(\mult_x_153/n43 ), .S(\mult_x_153/n45 ) );
  CMPE42D1BWP \mult_x_153/U31  ( .A(\mult_x_153/n149 ), .B(\mult_x_153/n127 ), 
        .C(\mult_x_153/n42 ), .CIX(\mult_x_153/n43 ), .D(\mult_x_153/n46 ), 
        .CO(\mult_x_153/n39 ), .COX(\mult_x_153/n38 ), .S(\mult_x_153/n40 ) );
  CMPE42D1BWP \mult_x_153/U29  ( .A(\mult_x_153/n137 ), .B(\mult_x_153/n37 ), 
        .C(\mult_x_153/n126 ), .CIX(\mult_x_153/n38 ), .D(\mult_x_153/n41 ), 
        .CO(\mult_x_153/n34 ), .COX(\mult_x_153/n33 ), .S(\mult_x_153/n35 ) );
  CMPE42D1BWP \mult_x_153/U28  ( .A(\mult_x_153/n117 ), .B(n6072), .C(
        \mult_x_153/n125 ), .CIX(\mult_x_153/n33 ), .D(\mult_x_153/n136 ), 
        .CO(\mult_x_153/n31 ), .COX(\mult_x_153/n30 ), .S(\mult_x_153/n32 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U55  ( .A1(\C1/Z_0 ), .A2(\C3/Z_0 ), .Z(
        \DP_OP_487J11_125_9213/n56 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U54  ( .A1(\C1/Z_0 ), .A2(\C3/Z_1 ), .Z(
        \DP_OP_487J11_125_9213/n55 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U53  ( .A1(\C1/Z_0 ), .A2(\C3/Z_2 ), .Z(
        \DP_OP_487J11_125_9213/n54 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U52  ( .A1(\C1/Z_0 ), .A2(\C3/Z_3 ), .Z(
        \DP_OP_487J11_125_9213/n53 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U51  ( .A1(\C1/Z_0 ), .A2(\C3/Z_4 ), .Z(
        \DP_OP_487J11_125_9213/n52 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U50  ( .A1(\C1/Z_0 ), .A2(\C3/Z_5 ), .Z(
        \DP_OP_487J11_125_9213/n51 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U49  ( .A1(\C1/Z_0 ), .A2(\C3/Z_6 ), .Z(
        \DP_OP_487J11_125_9213/n50 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U48  ( .A1(\C1/Z_0 ), .A2(\C3/Z_7 ), .Z(
        \DP_OP_487J11_125_9213/n49 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U47  ( .A1(\C1/Z_0 ), .A2(\C3/Z_8 ), .Z(
        \DP_OP_487J11_125_9213/n48 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U46  ( .A1(\C1/Z_0 ), .A2(\C3/Z_9 ), .Z(
        \DP_OP_487J11_125_9213/n47 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U45  ( .A1(\C1/Z_0 ), .A2(\C3/Z_10 ), .Z(
        \DP_OP_487J11_125_9213/n46 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U44  ( .A1(\C1/Z_0 ), .A2(\C3/Z_11 ), .Z(
        \DP_OP_487J11_125_9213/n45 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U43  ( .A1(\C1/Z_0 ), .A2(\C3/Z_12 ), .Z(
        \DP_OP_487J11_125_9213/n44 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U42  ( .A1(\C1/Z_0 ), .A2(\C3/Z_13 ), .Z(
        \DP_OP_487J11_125_9213/n43 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U41  ( .A1(\C1/Z_0 ), .A2(\C3/Z_14 ), .Z(
        \DP_OP_487J11_125_9213/n42 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U39  ( .A1(\C1/Z_0 ), .A2(\C3/Z_16 ), .Z(
        \DP_OP_487J11_125_9213/n40 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U38  ( .A1(\C1/Z_0 ), .A2(\C3/Z_17 ), .Z(
        \DP_OP_487J11_125_9213/n39 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U37  ( .A1(\C1/Z_0 ), .A2(\C3/Z_18 ), .Z(
        \DP_OP_487J11_125_9213/n38 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U36  ( .A1(\C1/Z_0 ), .A2(\C3/Z_19 ), .Z(
        \DP_OP_487J11_125_9213/n37 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U34  ( .A1(\C1/Z_0 ), .A2(\C3/Z_21 ), .Z(
        \DP_OP_487J11_125_9213/n35 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U33  ( .A1(\C1/Z_0 ), .A2(\C3/Z_22 ), .Z(
        \DP_OP_487J11_125_9213/n34 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U32  ( .A1(\C1/Z_0 ), .A2(\C3/Z_23 ), .Z(
        \DP_OP_487J11_125_9213/n33 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U31  ( .A1(\C1/Z_0 ), .A2(\C3/Z_24 ), .Z(
        \DP_OP_487J11_125_9213/n32 ) );
  XOR2D1BWP \DP_OP_487J11_125_9213/U30  ( .A1(\C1/Z_0 ), .A2(\C3/Z_25 ), .Z(
        \DP_OP_487J11_125_9213/n31 ) );
  FA1D0BWP \DP_OP_487J11_125_9213/U11  ( .A(\DP_OP_487J11_125_9213/n40 ), .B(
        \C2/Z_16 ), .CI(\DP_OP_487J11_125_9213/n11 ), .CO(
        \DP_OP_487J11_125_9213/n10 ), .S(N1473) );
  FA1D0BWP \DP_OP_487J11_125_9213/U10  ( .A(\DP_OP_487J11_125_9213/n39 ), .B(
        \C2/Z_17 ), .CI(\DP_OP_487J11_125_9213/n10 ), .CO(
        \DP_OP_487J11_125_9213/n9 ), .S(N1474) );
  FA1D0BWP \DP_OP_487J11_125_9213/U9  ( .A(\DP_OP_487J11_125_9213/n38 ), .B(
        \C2/Z_18 ), .CI(\DP_OP_487J11_125_9213/n9 ), .CO(
        \DP_OP_487J11_125_9213/n8 ), .S(N1475) );
  FA1D0BWP \DP_OP_487J11_125_9213/U8  ( .A(\DP_OP_487J11_125_9213/n37 ), .B(
        \C2/Z_19 ), .CI(\DP_OP_487J11_125_9213/n8 ), .CO(
        \DP_OP_487J11_125_9213/n7 ), .S(N1476) );
  FA1D0BWP \DP_OP_487J11_125_9213/U7  ( .A(\DP_OP_487J11_125_9213/n36 ), .B(
        \C2/Z_20 ), .CI(\DP_OP_487J11_125_9213/n7 ), .CO(
        \DP_OP_487J11_125_9213/n6 ), .S(N1477) );
  FA1D0BWP \DP_OP_487J11_125_9213/U6  ( .A(\DP_OP_487J11_125_9213/n35 ), .B(
        \C2/Z_21 ), .CI(\DP_OP_487J11_125_9213/n6 ), .CO(
        \DP_OP_487J11_125_9213/n5 ), .S(N1478) );
  FA1D0BWP \DP_OP_487J11_125_9213/U5  ( .A(\DP_OP_487J11_125_9213/n34 ), .B(
        \C2/Z_22 ), .CI(\DP_OP_487J11_125_9213/n5 ), .CO(
        \DP_OP_487J11_125_9213/n4 ), .S(N1479) );
  FA1D0BWP \DP_OP_487J11_125_9213/U4  ( .A(\DP_OP_487J11_125_9213/n33 ), .B(
        \C2/Z_23 ), .CI(\DP_OP_487J11_125_9213/n4 ), .CO(
        \DP_OP_487J11_125_9213/n3 ), .S(N1480) );
  FA1D0BWP \DP_OP_487J11_125_9213/U3  ( .A(\DP_OP_487J11_125_9213/n32 ), .B(
        \C2/Z_24 ), .CI(\DP_OP_487J11_125_9213/n3 ), .CO(
        \DP_OP_487J11_125_9213/n2 ), .S(N1481) );
  FA1D0BWP \DP_OP_487J11_125_9213/U2  ( .A(\DP_OP_487J11_125_9213/n31 ), .B(
        \C2/Z_25 ), .CI(\DP_OP_487J11_125_9213/n2 ), .CO(
        \DP_OP_487J11_125_9213/n1 ), .S(N1482) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U54  ( .A1(n4612), .A2(n4576), .Z(
        \DP_OP_493J11_130_7648/n55 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U53  ( .A1(n4612), .A2(n4577), .Z(
        \DP_OP_493J11_130_7648/n54 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U52  ( .A1(n4612), .A2(n4578), .Z(
        \DP_OP_493J11_130_7648/n53 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U51  ( .A1(n4612), .A2(n4579), .Z(
        \DP_OP_493J11_130_7648/n52 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U50  ( .A1(n4612), .A2(n4580), .Z(
        \DP_OP_493J11_130_7648/n51 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U49  ( .A1(n4612), .A2(n4581), .Z(
        \DP_OP_493J11_130_7648/n50 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U48  ( .A1(n4612), .A2(n4582), .Z(
        \DP_OP_493J11_130_7648/n49 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U47  ( .A1(n4612), .A2(n4583), .Z(
        \DP_OP_493J11_130_7648/n48 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U46  ( .A1(n4612), .A2(n4584), .Z(
        \DP_OP_493J11_130_7648/n47 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U45  ( .A1(n4612), .A2(n4585), .Z(
        \DP_OP_493J11_130_7648/n46 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U44  ( .A1(n4612), .A2(n4586), .Z(
        \DP_OP_493J11_130_7648/n45 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U43  ( .A1(n4612), .A2(n4587), .Z(
        \DP_OP_493J11_130_7648/n44 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U42  ( .A1(n4612), .A2(n4588), .Z(
        \DP_OP_493J11_130_7648/n43 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U41  ( .A1(n4612), .A2(n4589), .Z(
        \DP_OP_493J11_130_7648/n42 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U40  ( .A1(n4612), .A2(n4590), .Z(
        \DP_OP_493J11_130_7648/n41 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U39  ( .A1(n4612), .A2(n4591), .Z(
        \DP_OP_493J11_130_7648/n40 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U38  ( .A1(n4612), .A2(n4592), .Z(
        \DP_OP_493J11_130_7648/n39 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U37  ( .A1(n4612), .A2(n4593), .Z(
        \DP_OP_493J11_130_7648/n38 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U36  ( .A1(n4612), .A2(n4594), .Z(
        \DP_OP_493J11_130_7648/n37 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U35  ( .A1(n4612), .A2(n4595), .Z(
        \DP_OP_493J11_130_7648/n36 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U34  ( .A1(n4612), .A2(n4596), .Z(
        \DP_OP_493J11_130_7648/n35 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U33  ( .A1(n4612), .A2(n4597), .Z(
        \DP_OP_493J11_130_7648/n34 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U32  ( .A1(n4612), .A2(n4598), .Z(
        \DP_OP_493J11_130_7648/n33 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U31  ( .A1(n4612), .A2(n4599), .Z(
        \DP_OP_493J11_130_7648/n32 ) );
  XOR2D1BWP \DP_OP_493J11_130_7648/U30  ( .A1(n4612), .A2(n4600), .Z(
        \DP_OP_493J11_130_7648/n31 ) );
  FA1D0BWP \DP_OP_493J11_130_7648/U12  ( .A(\DP_OP_493J11_130_7648/n41 ), .B(
        n4601), .CI(\DP_OP_493J11_130_7648/n12 ), .CO(
        \DP_OP_493J11_130_7648/n11 ), .S(\alu/N328 ) );
  FA1D0BWP \DP_OP_493J11_130_7648/U11  ( .A(\DP_OP_493J11_130_7648/n40 ), .B(
        n4602), .CI(\DP_OP_493J11_130_7648/n11 ), .CO(
        \DP_OP_493J11_130_7648/n10 ), .S(\alu/N329 ) );
  FA1D0BWP \DP_OP_493J11_130_7648/U10  ( .A(\DP_OP_493J11_130_7648/n39 ), .B(
        n4603), .CI(\DP_OP_493J11_130_7648/n10 ), .CO(
        \DP_OP_493J11_130_7648/n9 ), .S(\alu/N330 ) );
  FA1D0BWP \DP_OP_493J11_130_7648/U9  ( .A(\DP_OP_493J11_130_7648/n38 ), .B(
        n4604), .CI(\DP_OP_493J11_130_7648/n9 ), .CO(
        \DP_OP_493J11_130_7648/n8 ), .S(\alu/N331 ) );
  FA1D0BWP \DP_OP_493J11_130_7648/U8  ( .A(\DP_OP_493J11_130_7648/n37 ), .B(
        n4605), .CI(\DP_OP_493J11_130_7648/n8 ), .CO(
        \DP_OP_493J11_130_7648/n7 ), .S(\alu/N332 ) );
  FA1D0BWP \DP_OP_493J11_130_7648/U7  ( .A(\DP_OP_493J11_130_7648/n36 ), .B(
        n4606), .CI(\DP_OP_493J11_130_7648/n7 ), .CO(
        \DP_OP_493J11_130_7648/n6 ), .S(\alu/N333 ) );
  FA1D0BWP \DP_OP_493J11_130_7648/U6  ( .A(\DP_OP_493J11_130_7648/n35 ), .B(
        n4607), .CI(\DP_OP_493J11_130_7648/n6 ), .CO(
        \DP_OP_493J11_130_7648/n5 ), .S(\alu/N334 ) );
  FA1D0BWP \DP_OP_493J11_130_7648/U5  ( .A(\DP_OP_493J11_130_7648/n34 ), .B(
        n4608), .CI(\DP_OP_493J11_130_7648/n5 ), .CO(
        \DP_OP_493J11_130_7648/n4 ), .S(\alu/N335 ) );
  FA1D0BWP \DP_OP_493J11_130_7648/U4  ( .A(\DP_OP_493J11_130_7648/n33 ), .B(
        n4609), .CI(\DP_OP_493J11_130_7648/n4 ), .CO(
        \DP_OP_493J11_130_7648/n3 ), .S(\alu/N336 ) );
  FA1D0BWP \DP_OP_493J11_130_7648/U3  ( .A(\DP_OP_493J11_130_7648/n32 ), .B(
        n4610), .CI(\DP_OP_493J11_130_7648/n3 ), .CO(
        \DP_OP_493J11_130_7648/n2 ), .S(\alu/N337 ) );
  FA1D0BWP \DP_OP_493J11_130_7648/U2  ( .A(\DP_OP_493J11_130_7648/n31 ), .B(
        n4611), .CI(\DP_OP_493J11_130_7648/n2 ), .CO(
        \DP_OP_493J11_130_7648/n1 ), .S(\alu/N338 ) );
  FA1D0BWP \intadd_33/U11  ( .A(\mult_x_153/n78 ), .B(\mult_x_153/n73 ), .CI(
        \intadd_33/CI ), .CO(\intadd_33/n10 ), .S(\intadd_33/SUM[0] ) );
  FA1D0BWP \intadd_33/U10  ( .A(\mult_x_153/n72 ), .B(\mult_x_153/n66 ), .CI(
        \intadd_33/n10 ), .CO(\intadd_33/n9 ), .S(\intadd_33/SUM[1] ) );
  FA1D0BWP \intadd_33/U9  ( .A(\mult_x_153/n58 ), .B(\mult_x_153/n65 ), .CI(
        \intadd_33/n9 ), .CO(\intadd_33/n8 ), .S(\intadd_33/SUM[2] ) );
  FA1D0BWP \intadd_33/U8  ( .A(\mult_x_153/n52 ), .B(\mult_x_153/n57 ), .CI(
        \intadd_33/n8 ), .CO(\intadd_33/n7 ), .S(\intadd_33/SUM[3] ) );
  FA1D0BWP \intadd_33/U7  ( .A(\mult_x_153/n45 ), .B(\mult_x_153/n51 ), .CI(
        \intadd_33/n7 ), .CO(\intadd_33/n6 ), .S(\intadd_33/SUM[4] ) );
  FA1D0BWP \intadd_33/U6  ( .A(\mult_x_153/n40 ), .B(\mult_x_153/n44 ), .CI(
        \intadd_33/n6 ), .CO(\intadd_33/n5 ), .S(\intadd_33/SUM[5] ) );
  FA1D0BWP \intadd_33/U5  ( .A(\mult_x_153/n35 ), .B(\mult_x_153/n39 ), .CI(
        \intadd_33/n5 ), .CO(\intadd_33/n4 ), .S(\intadd_33/SUM[6] ) );
  FA1D0BWP \intadd_33/U4  ( .A(\mult_x_153/n32 ), .B(\mult_x_153/n34 ), .CI(
        \intadd_33/n4 ), .CO(\intadd_33/n3 ), .S(\intadd_33/SUM[7] ) );
  FA1D0BWP \intadd_33/U3  ( .A(\mult_x_153/n31 ), .B(\intadd_33/B[8] ), .CI(
        \intadd_33/n3 ), .CO(\intadd_33/n2 ), .S(\intadd_33/SUM[8] ) );
  FA1D0BWP \intadd_33/U2  ( .A(\intadd_33/A[9] ), .B(\intadd_33/B[9] ), .CI(
        \intadd_33/n2 ), .CO(\intadd_33/n1 ), .S(\intadd_33/SUM[9] ) );
  FA1D0BWP \intadd_34/U3  ( .A(\intadd_34/A[2] ), .B(scalarToLoad[13]), .CI(
        \intadd_34/n3 ), .CO(\intadd_34/n2 ), .S(\intadd_34/SUM[2] ) );
  FA1D0BWP \intadd_34/U2  ( .A(\intadd_34/A[3] ), .B(scalarToLoad[14]), .CI(
        \intadd_34/n2 ), .CO(\intadd_34/n1 ), .S(\intadd_34/SUM[3] ) );
  FA1D0BWP \intadd_35/U4  ( .A(\intadd_35/A[0] ), .B(\intadd_35/B[0] ), .CI(
        \intadd_35/CI ), .CO(\intadd_35/n3 ), .S(\intadd_35/SUM[0] ) );
  FA1D0BWP \intadd_35/U3  ( .A(\intadd_35/A[1] ), .B(\intadd_35/B[1] ), .CI(
        \intadd_35/n3 ), .CO(\intadd_35/n2 ), .S(\intadd_35/SUM[1] ) );
  FA1D0BWP \intadd_35/U2  ( .A(\intadd_35/A[2] ), .B(\intadd_35/B[2] ), .CI(
        \intadd_35/n2 ), .CO(\intadd_35/n1 ), .S(\intadd_35/SUM[2] ) );
  FA1D0BWP \intadd_36/U4  ( .A(op2[11]), .B(\intadd_36/B[0] ), .CI(
        \intadd_36/CI ), .CO(\intadd_36/n3 ), .S(\intadd_36/SUM[0] ) );
  FA1D0BWP \intadd_36/U3  ( .A(op2[12]), .B(\intadd_36/B[1] ), .CI(
        \intadd_36/n3 ), .CO(\intadd_36/n2 ), .S(\intadd_36/SUM[1] ) );
  FA1D0BWP \intadd_36/U2  ( .A(op2[13]), .B(\intadd_36/B[2] ), .CI(
        \intadd_36/n2 ), .CO(\intadd_36/n1 ), .S(\intadd_36/SUM[2] ) );
  DFQD4BWP \state_reg[1]  ( .D(N153), .CP(Clk1), .Q(state[1]) );
  DFQD4BWP \state_reg[3]  ( .D(N155), .CP(Clk1), .Q(state[3]) );
  LHD1BWP \scalarToLoad_reg[13]  ( .E(n4695), .D(N1823), .Q(scalarToLoad[13]), 
        .QN(n3655) );
  LHD1BWP \op1_reg[13]  ( .E(N4208), .D(N4189), .Q(op1[13]), .QN(n3653) );
  LHD1BWP \wrAddr_reg[1]  ( .E(N4211), .D(N4213), .Q(n3651), .QN(n138) );
  LHD1BWP \scalarToLoad_reg[14]  ( .E(n4695), .D(N1824), .Q(scalarToLoad[14]), 
        .QN(n3638) );
  LHD1BWP \wrAddr_reg[0]  ( .E(N4211), .D(N4212), .Q(\srf/N15 ), .QN(n3637) );
  LHD1BWP \scalarToLoad_reg[10]  ( .E(n4695), .D(N1820), .Q(scalarToLoad[10]), 
        .QN(n3615) );
  LHD1BWP \vectorToLoad_reg[9]  ( .E(N4215), .D(N4225), .QN(n119) );
  LHD1BWP \vectorToLoad_reg[8]  ( .E(N4215), .D(N4224), .QN(n120) );
  LHD1BWP \vectorToLoad_reg[7]  ( .E(N4215), .D(N4223), .QN(n121) );
  LHD1BWP \vectorToLoad_reg[6]  ( .E(N4215), .D(N4222), .QN(n122) );
  LHD1BWP \vectorToLoad_reg[5]  ( .E(N4215), .D(N4221), .QN(n123) );
  LHD1BWP \vectorToLoad_reg[4]  ( .E(N4215), .D(N4220), .QN(n124) );
  LHD1BWP \vectorToLoad_reg[3]  ( .E(N4215), .D(N4219), .QN(n125) );
  LHD1BWP \vectorToLoad_reg[2]  ( .E(N4215), .D(N4218), .QN(n126) );
  LHD1BWP \vectorToLoad_reg[1]  ( .E(N4215), .D(N4217), .QN(n127) );
  LHD1BWP \vectorToLoad_reg[15]  ( .E(N4215), .D(N4231), .QN(n113) );
  LHD1BWP \vectorToLoad_reg[14]  ( .E(N4215), .D(N4230), .QN(n114) );
  LHD1BWP \vectorToLoad_reg[13]  ( .E(N4215), .D(N4229), .QN(n115) );
  LHD1BWP \vectorToLoad_reg[12]  ( .E(N4215), .D(N4228), .QN(n116) );
  LHD1BWP \vectorToLoad_reg[11]  ( .E(N4215), .D(N4227), .QN(n117) );
  LHD1BWP \vectorToLoad_reg[10]  ( .E(N4215), .D(N4226), .QN(n118) );
  LHD1BWP \vectorToLoad_reg[0]  ( .E(N4215), .D(N4216), .QN(n128) );
  LND1BWP \instrIn_reg[5]  ( .D(DataIn[5]), .EN(n3020), .QN(n153) );
  LHCNQD1BWP flow_reg ( .E(n4696), .D(overflow), .CDN(n156), .Q(V) );
  LHD1BWP \op2_reg[15]  ( .E(N4208), .D(N4207), .Q(op2[15]) );
  LHQD1BWP \func_reg[1]  ( .E(n4616), .D(n4697), .Q(n1) );
  LHQD1BWP \op2_reg[9]  ( .E(N4208), .D(N4201), .Q(op2[9]) );
  LHQD1BWP \op2_reg[5]  ( .E(N4208), .D(N4197), .Q(op2[5]) );
  LHQD1BWP \op2_reg[8]  ( .E(N4208), .D(N4200), .Q(op2[8]) );
  LHQD1BWP \op2_reg[6]  ( .E(N4208), .D(N4198), .Q(op2[6]) );
  LHD1BWP \scalarToLoad_reg[12]  ( .E(n4695), .D(N1822), .Q(scalarToLoad[12])
         );
  LHD1BWP \scalarToLoad_reg[11]  ( .E(n4695), .D(N1821), .Q(scalarToLoad[11])
         );
  LHD1BWP \op2_reg[13]  ( .E(N4208), .D(N4205), .Q(op2[13]), .QN(n3561) );
  LHQD1BWP \op2_reg[7]  ( .E(N4208), .D(N4199), .Q(op2[7]) );
  LHQD1BWP \wrAddr_reg[2]  ( .E(N4211), .D(N4214), .Q(\srf/N17 ) );
  LNQD1BWP \instrIn_reg[12]  ( .D(DataIn[12]), .EN(n3020), .Q(code[0]) );
  CKXOR2D0BWP \DP_OP_493J11_130_7648/U55  ( .A1(n4612), .A2(n4575), .Z(
        \DP_OP_493J11_130_7648/n56 ) );
  DFQD2BWP \state_reg[0]  ( .D(N152), .CP(Clk1), .Q(n3564) );
  DFQD4BWP \state_reg[2]  ( .D(n4614), .CP(Clk1), .Q(n3562) );
  CKND4BWP U4952 ( .I(state[1]), .ZN(n3663) );
  MOAI22D0BWP U4953 ( .A1(n3678), .A2(n4743), .B1(n4742), .B2(n3678), .ZN(
        n4750) );
  MOAI22D0BWP U4954 ( .A1(n3678), .A2(n4723), .B1(n4722), .B2(n3678), .ZN(
        n4730) );
  MOAI22D0BWP U4955 ( .A1(n4739), .A2(n3652), .B1(n3652), .B2(n4737), .ZN(
        n4741) );
  MOAI22D0BWP U4956 ( .A1(n4719), .A2(n3652), .B1(n3652), .B2(n4717), .ZN(
        n4720) );
  MOAI22D0BWP U4957 ( .A1(n5572), .A2(n5568), .B1(n5567), .B2(n5572), .ZN(
        n5578) );
  MOAI22D0BWP U4958 ( .A1(n4820), .A2(n4819), .B1(n4818), .B2(n4817), .ZN(
        \mult_x_153/n159 ) );
  MOAI22D0BWP U4959 ( .A1(n4825), .A2(n5562), .B1(n4824), .B2(n5572), .ZN(
        \mult_x_153/n168 ) );
  MOAI22D0BWP U4960 ( .A1(n4557), .A2(n4553), .B1(instrIn[3]), .B2(n4552), 
        .ZN(\vrf/N12 ) );
  MOAI22D0BWP U4961 ( .A1(n4560), .A2(n4553), .B1(instrIn[4]), .B2(n4552), 
        .ZN(\vrf/N13 ) );
  MOAI22D0BWP U4962 ( .A1(n5576), .A2(n4823), .B1(n4822), .B2(n5557), .ZN(
        \mult_x_153/n166 ) );
  MOAI22D0BWP U4963 ( .A1(n4430), .A2(n4429), .B1(\alu/N336 ), .B2(n4451), 
        .ZN(n4431) );
  MOAI22D0BWP U4964 ( .A1(n4207), .A2(n3676), .B1(n4318), .B2(n4216), .ZN(
        \C3/Z_17 ) );
  XNR2D1BWP U4965 ( .A1(\C1/Z_0 ), .A2(n3269), .ZN(\DP_OP_487J11_125_9213/n36 ) );
  AOI22D1BWP U4966 ( .A1(n4194), .A2(n4300), .B1(n4193), .B2(n4298), .ZN(n3269) );
  MOAI22D0BWP U4967 ( .A1(n4267), .A2(n4176), .B1(n4274), .B2(n4194), .ZN(
        \C3/Z_24 ) );
  MOAI22D0BWP U4968 ( .A1(n4258), .A2(n4166), .B1(n4326), .B2(n4194), .ZN(
        \C3/Z_25 ) );
  MAOI222D1BWP U4969 ( .A(n4352), .B(n4362), .C(n4358), .ZN(n4875) );
  MAOI222D1BWP U4970 ( .A(\mult_x_153/n91 ), .B(\mult_x_153/n85 ), .C(n5603), 
        .ZN(n5796) );
  ND2D1BWP U4971 ( .A1(n3565), .A2(n3563), .ZN(n3610) );
  IND2D1BWP U4972 ( .A1(n3598), .B1(n3663), .ZN(n3606) );
  MOAI22D0BWP U4973 ( .A1(n4561), .A2(n4555), .B1(instrIn[8]), .B2(n4554), 
        .ZN(\vrf/N11 ) );
  NR2XD0BWP U4974 ( .A1(n6074), .A2(n4622), .ZN(n6081) );
  NR2XD0BWP U4975 ( .A1(n6078), .A2(n4622), .ZN(n6083) );
  CKBD3BWP U4976 ( .I(n6081), .Z(n3573) );
  CKBD3BWP U4977 ( .I(n6075), .Z(n3593) );
  CKBD3BWP U4978 ( .I(n6083), .Z(n3578) );
  CKBD3BWP U4979 ( .I(n6079), .Z(n3597) );
  CKBD3BWP U4980 ( .I(n3573), .Z(n3591) );
  CKBD3BWP U4981 ( .I(n3593), .Z(n3566) );
  CKBD3BWP U4982 ( .I(n3578), .Z(n3592) );
  CKBD3BWP U4983 ( .I(n3597), .Z(n3568) );
  MOAI22D0BWP U4984 ( .A1(n5561), .A2(n5569), .B1(n5556), .B2(n4855), .ZN(
        n4854) );
  MOAI22D0BWP U4985 ( .A1(n4832), .A2(n5615), .B1(n4852), .B2(n4851), .ZN(
        n4850) );
  MOAI22D0BWP U4986 ( .A1(n5651), .A2(n5680), .B1(n5675), .B2(n5666), .ZN(
        n5652) );
  MAOI222D1BWP U4987 ( .A(op1[9]), .B(op2[9]), .C(n4843), .ZN(n4842) );
  CKBD1BWP U4988 ( .I(state[3]), .Z(n3612) );
  NR3D0BWP U4989 ( .A1(n3708), .A2(n3562), .A3(n4394), .ZN(n3709) );
  INR2D1BWP U4990 ( .A1(n3563), .B1(n3608), .ZN(n3607) );
  ND2D1BWP U4991 ( .A1(n4572), .A2(n4394), .ZN(n4398) );
  ND2D1BWP U4992 ( .A1(n3612), .A2(n3598), .ZN(n3604) );
  NR2XD0BWP U4993 ( .A1(n5999), .A2(Reset), .ZN(n6034) );
  NR2XD0BWP U4994 ( .A1(n6000), .A2(n6001), .ZN(n4469) );
  NR2XD0BWP U4995 ( .A1(Reset), .A2(n6040), .ZN(n6062) );
  CKBD3BWP U4996 ( .I(n3596), .Z(n3570) );
  CKBD3BWP U4997 ( .I(n3594), .Z(n3572) );
  CKBD3BWP U4998 ( .I(n3595), .Z(n3567) );
  CKBD3BWP U4999 ( .I(n3599), .Z(n3575) );
  NR2XD0BWP U5000 ( .A1(n4997), .A2(n5252), .ZN(n5184) );
  NR2XD0BWP U5001 ( .A1(n4996), .A2(n5252), .ZN(n5186) );
  NR2XD0BWP U5002 ( .A1(n4995), .A2(n5252), .ZN(n5188) );
  MAOI222D1BWP U5003 ( .A(n5812), .B(n4668), .C(n4968), .ZN(n4969) );
  MAOI222D1BWP U5004 ( .A(cycles[1]), .B(result[1]), .C(n5253), .ZN(n4968) );
  NR2XD1BWP U5005 ( .A1(n4543), .A2(n5252), .ZN(n4549) );
  INVD1BWP U5006 ( .I(n4473), .ZN(n4550) );
  NR2XD1BWP U5007 ( .A1(n4400), .A2(n4471), .ZN(n4548) );
  ND2D1BWP U5008 ( .A1(n4534), .A2(n4547), .ZN(n4407) );
  INR2D1BWP U5009 ( .A1(n4408), .B1(n132), .ZN(n4627) );
  INVD1BWP U5010 ( .I(n4627), .ZN(n5509) );
  CKND6BWP U5011 ( .I(n3562), .ZN(n3563) );
  NR3D1BWP U5012 ( .A1(n3782), .A2(n3563), .A3(n3664), .ZN(WR) );
  NR2XD0BWP U5013 ( .A1(n3783), .A2(n3782), .ZN(n4696) );
  INR2D1BWP U5014 ( .A1(\srf/N59 ), .B1(n6062), .ZN(\vrf/N296 ) );
  CKBD4BWP U5015 ( .I(\vrf/N296 ), .Z(n3590) );
  INR2D1BWP U5016 ( .A1(\srf/N58 ), .B1(n6062), .ZN(\vrf/N293 ) );
  CKBD4BWP U5017 ( .I(\vrf/N293 ), .Z(n3588) );
  INR2D1BWP U5018 ( .A1(\srf/N57 ), .B1(n6062), .ZN(\vrf/N290 ) );
  CKBD4BWP U5019 ( .I(\vrf/N290 ), .Z(n3589) );
  INR2D1BWP U5020 ( .A1(\srf/N56 ), .B1(n6062), .ZN(\vrf/N287 ) );
  CKBD4BWP U5021 ( .I(\vrf/N287 ), .Z(n3587) );
  INR2D1BWP U5022 ( .A1(\srf/N55 ), .B1(n6062), .ZN(\vrf/N284 ) );
  CKBD4BWP U5023 ( .I(\vrf/N284 ), .Z(n3586) );
  INR2D1BWP U5024 ( .A1(\srf/N54 ), .B1(n6062), .ZN(\vrf/N281 ) );
  CKBD4BWP U5025 ( .I(\vrf/N281 ), .Z(n3584) );
  INR2D1BWP U5026 ( .A1(\srf/N53 ), .B1(n6062), .ZN(\vrf/N278 ) );
  CKBD4BWP U5027 ( .I(\vrf/N278 ), .Z(n3585) );
  INR2D1BWP U5028 ( .A1(\srf/N36 ), .B1(n6062), .ZN(\vrf/N217 ) );
  CKBD4BWP U5029 ( .I(\vrf/N217 ), .Z(n3583) );
  MOAI22D0BWP U5030 ( .A1(n4979), .A2(n3614), .B1(n4061), .B2(
        nextInstrAddr[12]), .ZN(N4146) );
  NR2XD0BWP U5031 ( .A1(n4397), .A2(n4396), .ZN(n4630) );
  CKND2D0BWP U5032 ( .A1(n5715), .A2(n5717), .ZN(n3270) );
  NR3D0BWP U5033 ( .A1(n3270), .A2(n5712), .A3(n4445), .ZN(n5705) );
  NR4D0BWP U5034 ( .A1(\intadd_35/A[0] ), .A2(\intadd_35/A[2] ), .A3(n5695), 
        .A4(\intadd_35/A[1] ), .ZN(n3271) );
  ND3D0BWP U5035 ( .A1(\alu/N339 ), .A2(n4675), .A3(n3271), .ZN(n4460) );
  IND2D0BWP U5036 ( .A1(N1482), .B1(n4374), .ZN(n4376) );
  IAO21D0BWP U5037 ( .A1(n5796), .A2(n5797), .B(n5798), .ZN(n3272) );
  MUX2ND0BWP U5038 ( .I0(\mult_x_153/n84 ), .I1(n5799), .S(n3272), .ZN(n3273)
         );
  MOAI22D0BWP U5039 ( .A1(n5800), .A2(n3273), .B1(n5802), .B2(
        \intadd_33/SUM[0] ), .ZN(n3274) );
  AOI211D0BWP U5040 ( .A1(n4680), .A2(n4679), .B(n4054), .C(n4862), .ZN(n3275)
         );
  OAI22D0BWP U5041 ( .A1(n4679), .A2(n3912), .B1(n4680), .B2(n3913), .ZN(n3276) );
  AOI211D0BWP U5042 ( .A1(n3925), .A2(n3274), .B(n3275), .C(n3276), .ZN(n3277)
         );
  OAI21D0BWP U5043 ( .A1(n5748), .A2(n3901), .B(n3277), .ZN(result[0]) );
  IND2D0BWP U5044 ( .A1(n3732), .B1(n4392), .ZN(n3661) );
  AOI22D0BWP U5045 ( .A1(n5227), .A2(vectorData1[201]), .B1(n5187), .B2(
        vectorData1[233]), .ZN(n3278) );
  AOI22D0BWP U5046 ( .A1(n5232), .A2(vectorData1[153]), .B1(n5185), .B2(
        vectorData1[89]), .ZN(n3279) );
  ND4D0BWP U5047 ( .A1(n5080), .A2(n5081), .A3(n5082), .A4(n5083), .ZN(n3280)
         );
  AOI21D0BWP U5048 ( .A1(n5229), .A2(vectorData1[249]), .B(n3280), .ZN(n3281)
         );
  ND4D0BWP U5049 ( .A1(n7590), .A2(n7589), .A3(n7588), .A4(n7587), .ZN(n3282)
         );
  ND4D0BWP U5050 ( .A1(n7334), .A2(n7333), .A3(n7332), .A4(n7331), .ZN(n3283)
         );
  AOI22D0BWP U5051 ( .A1(n5231), .A2(n3282), .B1(n5188), .B2(n3283), .ZN(n3284) );
  AN4D0BWP U5052 ( .A1(n3278), .A2(n3279), .A3(n3281), .A4(n3284), .Z(n3285)
         );
  AOI22D0BWP U5053 ( .A1(n8278), .A2(\srf/regTable[0][9] ), .B1(n8280), .B2(
        \srf/regTable[2][9] ), .ZN(n3286) );
  AOI22D0BWP U5054 ( .A1(n8284), .A2(\srf/regTable[3][9] ), .B1(n8282), .B2(
        \srf/regTable[1][9] ), .ZN(n3287) );
  AOI22D0BWP U5055 ( .A1(n8285), .A2(\srf/regTable[4][9] ), .B1(n8286), .B2(
        \srf/regTable[6][9] ), .ZN(n3288) );
  AOI22D0BWP U5056 ( .A1(n8288), .A2(\srf/regTable[7][9] ), .B1(n8287), .B2(
        \srf/regTable[5][9] ), .ZN(n3289) );
  ND4D0BWP U5057 ( .A1(n3286), .A2(n3287), .A3(n3288), .A4(n3289), .ZN(n3290)
         );
  AOI22D0BWP U5058 ( .A1(n3572), .A2(\vrf/regTable[2][9] ), .B1(n3581), .B2(
        \vrf/regTable[0][9] ), .ZN(n3291) );
  AOI22D0BWP U5059 ( .A1(n3579), .A2(\vrf/regTable[1][9] ), .B1(n3575), .B2(
        \vrf/regTable[3][9] ), .ZN(n3292) );
  AOI22D0BWP U5060 ( .A1(n3570), .A2(\vrf/regTable[6][9] ), .B1(n3574), .B2(
        \vrf/regTable[4][9] ), .ZN(n3293) );
  AOI22D0BWP U5061 ( .A1(n3576), .A2(\vrf/regTable[5][9] ), .B1(n3567), .B2(
        \vrf/regTable[7][9] ), .ZN(n3294) );
  ND4D0BWP U5062 ( .A1(n3291), .A2(n3292), .A3(n3293), .A4(n3294), .ZN(n3295)
         );
  AOI22D0BWP U5063 ( .A1(n4073), .A2(n3290), .B1(n4072), .B2(n3295), .ZN(n3296) );
  CKND2D0BWP U5064 ( .A1(n4071), .A2(Addr[9]), .ZN(n3297) );
  OAI211D0BWP U5065 ( .A1(n4070), .A2(n3285), .B(n3296), .C(n3297), .ZN(N4185)
         );
  AOI22D0BWP U5066 ( .A1(result[10]), .A2(n4975), .B1(n4699), .B2(n4976), .ZN(
        n3298) );
  MOAI22D0BWP U5067 ( .A1(n3614), .A2(n3298), .B1(n4061), .B2(
        nextInstrAddr[10]), .ZN(N4144) );
  IND2D0BWP U5068 ( .A1(n3799), .B1(n3800), .ZN(n3889) );
  CKND0BWP U5069 ( .I(n4153), .ZN(n3299) );
  AOI222D0BWP U5070 ( .A1(n3299), .A2(n4636), .B1(n4341), .B2(N1476), .C1(
        N1483), .C2(N1477), .ZN(n3300) );
  IOA21D0BWP U5071 ( .A1(n4373), .A2(n4152), .B(n3300), .ZN(n4896) );
  MUX2ND0BWP U5072 ( .I0(n5770), .I1(n5777), .S(n5778), .ZN(n3301) );
  MUX2ND0BWP U5073 ( .I0(n3301), .I1(n5770), .S(n5775), .ZN(n3302) );
  CKND0BWP U5074 ( .I(n5790), .ZN(n3303) );
  AOI211D0BWP U5075 ( .A1(n5774), .A2(n5773), .B(n5772), .C(n5771), .ZN(n3304)
         );
  XNR2D0BWP U5076 ( .A1(n3301), .A2(n3304), .ZN(n3305) );
  AOI22D0BWP U5077 ( .A1(n3301), .A2(n5786), .B1(n3303), .B2(n3305), .ZN(n3306) );
  OAI211D0BWP U5078 ( .A1(n5776), .A2(n3302), .B(n4656), .C(n3306), .ZN(n3307)
         );
  AOI22D0BWP U5079 ( .A1(op1[12]), .A2(n4672), .B1(n4689), .B2(n3307), .ZN(
        n3308) );
  AOI22D0BWP U5080 ( .A1(op2[4]), .A2(n4671), .B1(n4690), .B2(\alu/N1016 ), 
        .ZN(n3309) );
  OAI211D0BWP U5081 ( .A1(n5686), .A2(n5685), .B(n5804), .C(n5687), .ZN(n3310)
         );
  OAI21D0BWP U5082 ( .A1(n4691), .A2(n4692), .B(n3310), .ZN(n3311) );
  ND3D0BWP U5083 ( .A1(n3308), .A2(n3309), .A3(n3311), .ZN(result[12]) );
  AOI22D0BWP U5084 ( .A1(n5232), .A2(vectorData2[151]), .B1(n5227), .B2(
        vectorData2[199]), .ZN(n3312) );
  AO22D0BWP U5085 ( .A1(n5233), .A2(vectorData2[183]), .B1(n5228), .B2(
        vectorData2[215]), .Z(n3313) );
  AOI22D0BWP U5086 ( .A1(n5185), .A2(vectorData2[87]), .B1(n3601), .B2(
        vectorData2[39]), .ZN(n3314) );
  AOI22D0BWP U5087 ( .A1(n5226), .A2(vectorData2[135]), .B1(n5184), .B2(
        vectorData2[23]), .ZN(n3315) );
  AOI22D0BWP U5088 ( .A1(n5229), .A2(vectorData2[247]), .B1(n5230), .B2(
        vectorData2[167]), .ZN(n3316) );
  AOI22D0BWP U5089 ( .A1(n5186), .A2(vectorData2[71]), .B1(n5231), .B2(
        vectorData2[119]), .ZN(n3317) );
  ND4D0BWP U5090 ( .A1(n3314), .A2(n3315), .A3(n3316), .A4(n3317), .ZN(n3318)
         );
  AOI211D0BWP U5091 ( .A1(n5187), .A2(vectorData2[231]), .B(n3313), .C(n3318), 
        .ZN(n3319) );
  AOI22D0BWP U5092 ( .A1(n3671), .A2(vectorData2[103]), .B1(n5188), .B2(
        vectorData2[55]), .ZN(n3320) );
  AOI31D0BWP U5093 ( .A1(n3312), .A2(n3319), .A3(n3320), .B(n3661), .ZN(n3321)
         );
  AOI211D0BWP U5094 ( .A1(n4681), .A2(vectorData2[7]), .B(n5200), .C(n3321), 
        .ZN(n3322) );
  CKND2D0BWP U5095 ( .A1(n4688), .A2(scalarData2[7]), .ZN(n3323) );
  OAI211D0BWP U5096 ( .A1(n3883), .A2(n4559), .B(n3322), .C(n3323), .ZN(N4199)
         );
  AOI222D0BWP U5097 ( .A1(n5230), .A2(vectorData1[170]), .B1(n5233), .B2(
        vectorData1[186]), .C1(n3601), .C2(vectorData1[42]), .ZN(n3324) );
  IOA21D0BWP U5098 ( .A1(n5232), .A2(vectorData1[154]), .B(n3324), .ZN(n3325)
         );
  AOI211D0BWP U5099 ( .A1(vectorData1[90]), .A2(n5185), .B(n5088), .C(n3325), 
        .ZN(n3326) );
  AOI22D0BWP U5100 ( .A1(n8278), .A2(\srf/regTable[0][10] ), .B1(n8280), .B2(
        \srf/regTable[2][10] ), .ZN(n3327) );
  AOI22D0BWP U5101 ( .A1(n8284), .A2(\srf/regTable[3][10] ), .B1(n8282), .B2(
        \srf/regTable[1][10] ), .ZN(n3328) );
  AOI22D0BWP U5102 ( .A1(n8285), .A2(\srf/regTable[4][10] ), .B1(n8286), .B2(
        \srf/regTable[6][10] ), .ZN(n3329) );
  AOI22D0BWP U5103 ( .A1(n8288), .A2(\srf/regTable[7][10] ), .B1(n8287), .B2(
        \srf/regTable[5][10] ), .ZN(n3330) );
  ND4D0BWP U5104 ( .A1(n3327), .A2(n3328), .A3(n3329), .A4(n3330), .ZN(n3331)
         );
  AOI22D0BWP U5105 ( .A1(n3581), .A2(\vrf/regTable[0][10] ), .B1(n3572), .B2(
        \vrf/regTable[2][10] ), .ZN(n3332) );
  AOI22D0BWP U5106 ( .A1(n3579), .A2(\vrf/regTable[1][10] ), .B1(n3575), .B2(
        \vrf/regTable[3][10] ), .ZN(n3333) );
  AOI22D0BWP U5107 ( .A1(n3574), .A2(\vrf/regTable[4][10] ), .B1(n3570), .B2(
        \vrf/regTable[6][10] ), .ZN(n3334) );
  AOI22D0BWP U5108 ( .A1(n3576), .A2(\vrf/regTable[5][10] ), .B1(n3567), .B2(
        \vrf/regTable[7][10] ), .ZN(n3335) );
  ND4D0BWP U5109 ( .A1(n3332), .A2(n3333), .A3(n3334), .A4(n3335), .ZN(n3336)
         );
  CKND0BWP U5110 ( .I(n3830), .ZN(n3337) );
  AOI222D0BWP U5111 ( .A1(n3331), .A2(n4073), .B1(n3336), .B2(n4072), .C1(
        n3337), .C2(Addr[10]), .ZN(n3338) );
  ND4D0BWP U5112 ( .A1(n7530), .A2(n7529), .A3(n7528), .A4(n7527), .ZN(n3339)
         );
  ND4D0BWP U5113 ( .A1(n7338), .A2(n7337), .A3(n7336), .A4(n7335), .ZN(n3340)
         );
  AOI22D0BWP U5114 ( .A1(n5213), .A2(n3339), .B1(n5188), .B2(n3340), .ZN(n3341) );
  AOI32D0BWP U5115 ( .A1(n3326), .A2(n3338), .A3(n3341), .B1(n4070), .B2(n3338), .ZN(N4186) );
  OAI21D0BWP U5116 ( .A1(cycles[4]), .A2(n4970), .B(n4972), .ZN(n3342) );
  MOAI22D0BWP U5117 ( .A1(n3614), .A2(n3342), .B1(n4061), .B2(nextInstrAddr[4]), .ZN(N4138) );
  CKMUX2D0BWP U5118 ( .I0(N1475), .I1(N1476), .S(n4355), .Z(n4124) );
  CKND0BWP U5119 ( .I(n4674), .ZN(n3343) );
  AOI222D0BWP U5120 ( .A1(n3890), .A2(n3343), .B1(n3890), .B2(n3889), .C1(
        n4645), .C2(n4674), .ZN(n4644) );
  OAI32D0BWP U5121 ( .A1(n4929), .A2(n4913), .A3(n4912), .B1(n4930), .B2(n4929), .ZN(n3344) );
  OAI21D0BWP U5122 ( .A1(n3344), .A2(n4927), .B(n4928), .ZN(n3345) );
  CKND0BWP U5123 ( .I(n4932), .ZN(n3346) );
  AOI32D0BWP U5124 ( .A1(n4931), .A2(n4940), .A3(n3345), .B1(n3346), .B2(n4940), .ZN(n4942) );
  IND2D0BWP U5125 ( .A1(n5816), .B1(n5294), .ZN(n4472) );
  IOA21D0BWP U5126 ( .A1(n5290), .A2(n5291), .B(n5292), .ZN(n5419) );
  AOI21D0BWP U5127 ( .A1(n5767), .A2(n5765), .B(n5771), .ZN(n3347) );
  NR2D0BWP U5128 ( .A1(n5769), .A2(n5776), .ZN(n3348) );
  AOI22D0BWP U5129 ( .A1(n5767), .A2(n5766), .B1(n5768), .B2(n3348), .ZN(n3349) );
  OAI211D0BWP U5130 ( .A1(n5790), .A2(n3347), .B(n4656), .C(n3349), .ZN(n3350)
         );
  AOI22D0BWP U5131 ( .A1(op1[11]), .A2(n4672), .B1(n4689), .B2(n3350), .ZN(
        n3351) );
  AOI22D0BWP U5132 ( .A1(op2[3]), .A2(n4671), .B1(n4690), .B2(\alu/N1015 ), 
        .ZN(n3352) );
  CKND2D0BWP U5133 ( .A1(n5803), .A2(n5684), .ZN(n3353) );
  OAI211D0BWP U5134 ( .A1(n5803), .A2(n5684), .B(n5804), .C(n3353), .ZN(n3354)
         );
  OAI21D0BWP U5135 ( .A1(n4691), .A2(n4692), .B(n3354), .ZN(n3355) );
  ND3D0BWP U5136 ( .A1(n3351), .A2(n3352), .A3(n3355), .ZN(result[11]) );
  AOI22D0BWP U5137 ( .A1(n5232), .A2(vectorData2[150]), .B1(n5185), .B2(
        vectorData2[86]), .ZN(n3356) );
  AO22D0BWP U5138 ( .A1(n5233), .A2(vectorData2[182]), .B1(n5188), .B2(
        vectorData2[54]), .Z(n3357) );
  AOI22D0BWP U5139 ( .A1(n5231), .A2(vectorData2[118]), .B1(n3601), .B2(
        vectorData2[38]), .ZN(n3358) );
  AOI22D0BWP U5140 ( .A1(n5227), .A2(vectorData2[198]), .B1(n5229), .B2(
        vectorData2[246]), .ZN(n3359) );
  AOI22D0BWP U5141 ( .A1(n5230), .A2(vectorData2[166]), .B1(n5226), .B2(
        vectorData2[134]), .ZN(n3360) );
  AOI22D0BWP U5142 ( .A1(n5228), .A2(vectorData2[214]), .B1(n5184), .B2(
        vectorData2[22]), .ZN(n3361) );
  ND4D0BWP U5143 ( .A1(n3358), .A2(n3359), .A3(n3360), .A4(n3361), .ZN(n3362)
         );
  AOI211D0BWP U5144 ( .A1(n3671), .A2(vectorData2[102]), .B(n3357), .C(n3362), 
        .ZN(n3363) );
  AOI22D0BWP U5145 ( .A1(n5186), .A2(vectorData2[70]), .B1(n5187), .B2(
        vectorData2[230]), .ZN(n3364) );
  AOI31D0BWP U5146 ( .A1(n3356), .A2(n3363), .A3(n3364), .B(n3661), .ZN(n3365)
         );
  AOI211D0BWP U5147 ( .A1(n4681), .A2(vectorData2[6]), .B(n5200), .C(n3365), 
        .ZN(n3366) );
  CKND2D0BWP U5148 ( .A1(n4688), .A2(scalarData2[6]), .ZN(n3367) );
  OAI211D0BWP U5149 ( .A1(n3883), .A2(n4556), .B(n3366), .C(n3367), .ZN(N4198)
         );
  MUX2ND0BWP U5150 ( .I0(n6011), .I1(result[3]), .S(n4969), .ZN(n3368) );
  MUX2ND0BWP U5151 ( .I0(cycles[3]), .I1(n3675), .S(n3368), .ZN(n3369) );
  MOAI22D0BWP U5152 ( .A1(n3614), .A2(n3369), .B1(n4061), .B2(nextInstrAddr[3]), .ZN(N4137) );
  CKND0BWP U5153 ( .I(n4449), .ZN(n3370) );
  AOI22D0BWP U5154 ( .A1(\alu/N336 ), .A2(\alu/N335 ), .B1(\alu/N334 ), .B2(
        n3370), .ZN(n3371) );
  AOI22D0BWP U5155 ( .A1(\alu/N339 ), .A2(\alu/N338 ), .B1(\alu/N336 ), .B2(
        n4450), .ZN(n3372) );
  MAOI22D0BWP U5156 ( .A1(n4453), .A2(n4454), .B1(n4448), .B2(n4447), .ZN(
        n3373) );
  OAI211D0BWP U5157 ( .A1(n4452), .A2(n3371), .B(n3372), .C(n3373), .ZN(n3374)
         );
  AOI21D0BWP U5158 ( .A1(\alu/N337 ), .A2(n4451), .B(n3374), .ZN(n4624) );
  CKND0BWP U5159 ( .I(\C1/Z_0 ), .ZN(n3375) );
  AOI222D0BWP U5160 ( .A1(n4273), .A2(n4280), .B1(n4302), .B2(n4279), .C1(
        n4242), .C2(n4306), .ZN(n3376) );
  AOI22D0BWP U5161 ( .A1(n4302), .A2(n4281), .B1(n4246), .B2(n4282), .ZN(n3377) );
  OAI22D0BWP U5162 ( .A1(\intadd_34/n1 ), .A2(n3376), .B1(n3676), .B2(n3377), 
        .ZN(n3378) );
  MUX2ND0BWP U5163 ( .I0(\C1/Z_0 ), .I1(n3375), .S(n3378), .ZN(n3379) );
  OA22D1BWP U5164 ( .A1(\intadd_34/CO ), .A2(n6004), .B1(n3676), .B2(n4240), 
        .Z(n3380) );
  CKND2D0BWP U5165 ( .A1(\DP_OP_487J11_125_9213/n13 ), .A2(
        \DP_OP_487J11_125_9213/n42 ), .ZN(n3381) );
  MAOI222D0BWP U5166 ( .A(n3379), .B(n3380), .C(n3381), .ZN(
        \DP_OP_487J11_125_9213/n11 ) );
  XNR3D0BWP U5167 ( .A1(n3380), .A2(n3379), .A3(n3381), .ZN(N1472) );
  IND2D0BWP U5168 ( .A1(n4894), .B1(n4895), .ZN(n4353) );
  AN4D0BWP U5169 ( .A1(n4907), .A2(n4905), .A3(n4871), .A4(n4869), .Z(n4955)
         );
  INR2D0BWP U5170 ( .A1(n5184), .B1(n3661), .ZN(n4685) );
  AOI22D0BWP U5171 ( .A1(n5802), .A2(\intadd_33/SUM[5] ), .B1(n5801), .B2(
        \intadd_33/SUM[4] ), .ZN(n3382) );
  CKND0BWP U5172 ( .I(n3925), .ZN(n3383) );
  AOI22D0BWP U5173 ( .A1(op2[5]), .A2(n4672), .B1(op1[5]), .B2(n4671), .ZN(
        n3384) );
  ND3D0BWP U5174 ( .A1(n4656), .A2(n5761), .A3(n5737), .ZN(n3385) );
  CKND0BWP U5175 ( .I(n5738), .ZN(n3386) );
  MUX4ND0BWP U5176 ( .I0(n5744), .I1(n3386), .I2(n5741), .I3(n5746), .S0(n5772), .S1(n5745), .ZN(n3387) );
  OAI22D0BWP U5177 ( .A1(n5736), .A2(n5754), .B1(n3385), .B2(n3387), .ZN(n3388) );
  MUX2ND0BWP U5178 ( .I0(n4853), .I1(n4852), .S(n4851), .ZN(n3389) );
  AOI22D0BWP U5179 ( .A1(n4689), .A2(n3388), .B1(n4690), .B2(n3389), .ZN(n3390) );
  OAI211D0BWP U5180 ( .A1(n3382), .A2(n3383), .B(n3384), .C(n3390), .ZN(
        result[5]) );
  AOI222D0BWP U5181 ( .A1(n5232), .A2(vectorData1[155]), .B1(n5226), .B2(
        vectorData1[139]), .C1(n3671), .C2(vectorData1[107]), .ZN(n3391) );
  IOA21D0BWP U5182 ( .A1(n5187), .A2(vectorData1[235]), .B(n3391), .ZN(n3392)
         );
  AOI211D0BWP U5183 ( .A1(vectorData1[251]), .A2(n5229), .B(n5093), .C(n3392), 
        .ZN(n3393) );
  AOI22D0BWP U5184 ( .A1(n8278), .A2(\srf/regTable[0][11] ), .B1(n8280), .B2(
        \srf/regTable[2][11] ), .ZN(n3394) );
  AOI22D0BWP U5185 ( .A1(n8284), .A2(\srf/regTable[3][11] ), .B1(n8282), .B2(
        \srf/regTable[1][11] ), .ZN(n3395) );
  AOI22D0BWP U5186 ( .A1(n8285), .A2(\srf/regTable[4][11] ), .B1(n8286), .B2(
        \srf/regTable[6][11] ), .ZN(n3396) );
  AOI22D0BWP U5187 ( .A1(n8288), .A2(\srf/regTable[7][11] ), .B1(n8287), .B2(
        \srf/regTable[5][11] ), .ZN(n3397) );
  ND4D0BWP U5188 ( .A1(n3394), .A2(n3395), .A3(n3396), .A4(n3397), .ZN(n3398)
         );
  AOI22D0BWP U5189 ( .A1(n3581), .A2(\vrf/regTable[0][11] ), .B1(n3572), .B2(
        \vrf/regTable[2][11] ), .ZN(n3399) );
  AOI22D0BWP U5190 ( .A1(n3579), .A2(\vrf/regTable[1][11] ), .B1(n3575), .B2(
        \vrf/regTable[3][11] ), .ZN(n3400) );
  AOI22D0BWP U5191 ( .A1(n3574), .A2(\vrf/regTable[4][11] ), .B1(n3570), .B2(
        \vrf/regTable[6][11] ), .ZN(n3401) );
  AOI22D0BWP U5192 ( .A1(n3576), .A2(\vrf/regTable[5][11] ), .B1(n3567), .B2(
        \vrf/regTable[7][11] ), .ZN(n3402) );
  ND4D0BWP U5193 ( .A1(n3399), .A2(n3400), .A3(n3401), .A4(n3402), .ZN(n3403)
         );
  CKND0BWP U5194 ( .I(n3830), .ZN(n3404) );
  AOI222D0BWP U5195 ( .A1(n3398), .A2(n4073), .B1(n3403), .B2(n4072), .C1(
        n3404), .C2(Addr[11]), .ZN(n3405) );
  ND4D0BWP U5196 ( .A1(n7598), .A2(n7597), .A3(n7596), .A4(n7595), .ZN(n3406)
         );
  ND4D0BWP U5197 ( .A1(n7406), .A2(n7405), .A3(n7404), .A4(n7403), .ZN(n3407)
         );
  AOI22D0BWP U5198 ( .A1(n5231), .A2(n3406), .B1(n5186), .B2(n3407), .ZN(n3408) );
  AOI32D0BWP U5199 ( .A1(n3393), .A2(n3405), .A3(n3408), .B1(n4070), .B2(n3405), .ZN(N4187) );
  MUX2ND0BWP U5200 ( .I0(result[2]), .I1(n4668), .S(n4968), .ZN(n3409) );
  MUX2ND0BWP U5201 ( .I0(cycles[2]), .I1(n5812), .S(n3409), .ZN(n3410) );
  MOAI22D0BWP U5202 ( .A1(n3614), .A2(n3410), .B1(n4061), .B2(nextInstrAddr[2]), .ZN(N4136) );
  MOAI22D0BWP U5203 ( .A1(n4797), .A2(n5554), .B1(n4796), .B2(n4795), .ZN(
        \mult_x_153/n133 ) );
  MOAI22D0BWP U5204 ( .A1(n4808), .A2(n4807), .B1(n4806), .B2(n4805), .ZN(
        \mult_x_153/n144 ) );
  AN2D0BWP U5205 ( .A1(\DP_OP_487J11_125_9213/n14 ), .A2(
        \DP_OP_487J11_125_9213/n43 ), .Z(\DP_OP_487J11_125_9213/n13 ) );
  AOI22D0BWP U5206 ( .A1(\alu/N339 ), .A2(\alu/N336 ), .B1(\alu/N334 ), .B2(
        n4450), .ZN(n3411) );
  CKND2D0BWP U5207 ( .A1(n4451), .A2(\alu/N335 ), .ZN(n3412) );
  OAI211D0BWP U5208 ( .A1(n4452), .A2(n4440), .B(n3411), .C(n3412), .ZN(n3413)
         );
  AOI21D0BWP U5209 ( .A1(n4453), .A2(n4427), .B(n3413), .ZN(n3414) );
  OAI31D0BWP U5210 ( .A1(\intadd_35/B[0] ), .A2(n4448), .A3(n4425), .B(n3414), 
        .ZN(n4446) );
  CKND0BWP U5211 ( .I(n4901), .ZN(n3415) );
  CKND0BWP U5212 ( .I(n4902), .ZN(n3416) );
  CKND2D0BWP U5213 ( .A1(n4871), .A2(n4870), .ZN(n3417) );
  OAI221D0BWP U5214 ( .A1(n4904), .A2(n4871), .B1(n4870), .B2(n4907), .C(n3417), .ZN(n3418) );
  CKND0BWP U5215 ( .I(n4899), .ZN(n3419) );
  OAI22D0BWP U5216 ( .A1(n3419), .A2(n4898), .B1(n4894), .B2(n4895), .ZN(n3420) );
  AOI221D0BWP U5217 ( .A1(n3419), .A2(n4898), .B1(n4895), .B2(n4894), .C(n3420), .ZN(n3421) );
  CKND0BWP U5218 ( .I(n4634), .ZN(n3422) );
  CKND0BWP U5219 ( .I(n4353), .ZN(n3423) );
  OAI22D0BWP U5220 ( .A1(n3422), .A2(n4896), .B1(n3423), .B2(n4354), .ZN(n3424) );
  AOI221D0BWP U5221 ( .A1(n3422), .A2(n4896), .B1(n4354), .B2(n3423), .C(n3424), .ZN(n3425) );
  IND4D0BWP U5222 ( .A1(n4868), .B1(n4892), .B2(n3421), .B3(n3425), .ZN(n3426)
         );
  AOI211D0BWP U5223 ( .A1(n4907), .A2(n4904), .B(n3418), .C(n3426), .ZN(n3427)
         );
  OAI221D0BWP U5224 ( .A1(n4902), .A2(n3415), .B1(n3416), .B2(n4901), .C(n3427), .ZN(n4888) );
  IND2D0BWP U5225 ( .A1(n4542), .B1(n3732), .ZN(n4572) );
  INR2D0BWP U5226 ( .A1(n5188), .B1(n3661), .ZN(n4686) );
  NR2D0BWP U5227 ( .A1(n4691), .A2(n4692), .ZN(n3428) );
  CKND0BWP U5228 ( .I(n5804), .ZN(n3429) );
  AOI211D0BWP U5229 ( .A1(n5688), .A2(n5687), .B(n5690), .C(n3429), .ZN(n3430)
         );
  CKND2D0BWP U5230 ( .A1(n5777), .A2(n5778), .ZN(n3431) );
  MUX2ND0BWP U5231 ( .I0(n5779), .I1(n5780), .S(n3431), .ZN(n3432) );
  NR2D0BWP U5232 ( .A1(n5776), .A2(n5787), .ZN(n3433) );
  CKND0BWP U5233 ( .I(n5781), .ZN(n3434) );
  AOI222D0BWP U5234 ( .A1(n3432), .A2(n3433), .B1(n3432), .B2(n5786), .C1(
        n3433), .C2(n3434), .ZN(n3435) );
  CKND2D0BWP U5235 ( .A1(n4656), .A2(n3435), .ZN(n3436) );
  AOI22D0BWP U5236 ( .A1(op1[13]), .A2(n4672), .B1(n4689), .B2(n3436), .ZN(
        n3437) );
  MUX2ND0BWP U5237 ( .I0(n4839), .I1(n4838), .S(n4837), .ZN(n3438) );
  AOI22D0BWP U5238 ( .A1(op2[5]), .A2(n4671), .B1(n4690), .B2(n3438), .ZN(
        n3439) );
  OAI211D0BWP U5239 ( .A1(n3428), .A2(n3430), .B(n3437), .C(n3439), .ZN(
        result[13]) );
  MUX2ND0BWP U5240 ( .I0(n4643), .I1(result[1]), .S(n5253), .ZN(n3440) );
  MUX2ND0BWP U5241 ( .I0(cycles[1]), .I1(n5417), .S(n3440), .ZN(n3441) );
  MOAI22D0BWP U5242 ( .A1(n3614), .A2(n3441), .B1(n4061), .B2(nextInstrAddr[1]), .ZN(N4135) );
  AN2D0BWP U5243 ( .A1(\DP_OP_493J11_130_7648/n16 ), .A2(
        \DP_OP_493J11_130_7648/n45 ), .Z(\DP_OP_493J11_130_7648/n15 ) );
  AN2D0BWP U5244 ( .A1(\DP_OP_493J11_130_7648/n20 ), .A2(
        \DP_OP_493J11_130_7648/n49 ), .Z(\DP_OP_493J11_130_7648/n19 ) );
  AN2D0BWP U5245 ( .A1(\DP_OP_493J11_130_7648/n24 ), .A2(
        \DP_OP_493J11_130_7648/n53 ), .Z(\DP_OP_493J11_130_7648/n23 ) );
  AN2D0BWP U5246 ( .A1(\DP_OP_487J11_125_9213/n17 ), .A2(
        \DP_OP_487J11_125_9213/n46 ), .Z(\DP_OP_487J11_125_9213/n16 ) );
  AN2D0BWP U5247 ( .A1(\DP_OP_487J11_125_9213/n23 ), .A2(
        \DP_OP_487J11_125_9213/n52 ), .Z(\DP_OP_487J11_125_9213/n22 ) );
  MOAI22D0BWP U5248 ( .A1(n4816), .A2(n4819), .B1(n4815), .B2(n4814), .ZN(
        \mult_x_153/n158 ) );
  INR2D0BWP U5249 ( .A1(n5703), .B1(n3885), .ZN(n3870) );
  IND2D0BWP U5250 ( .A1(n4887), .B1(n4866), .ZN(n4369) );
  CKND0BWP U5251 ( .I(n5718), .ZN(n3442) );
  CKND0BWP U5252 ( .I(n5720), .ZN(n3443) );
  AOI32D0BWP U5253 ( .A1(n5721), .A2(n3442), .A3(n3443), .B1(n4446), .B2(n3442), .ZN(n5755) );
  IND2D0BWP U5254 ( .A1(n4903), .B1(n4634), .ZN(n4156) );
  CKND0BWP U5255 ( .I(result[4]), .ZN(n3444) );
  OAI21D0BWP U5256 ( .A1(n4971), .A2(n3444), .B(n4972), .ZN(n4973) );
  AOI22D0BWP U5257 ( .A1(n5802), .A2(\intadd_33/SUM[9] ), .B1(n5801), .B2(
        \intadd_33/SUM[8] ), .ZN(n3445) );
  CKND0BWP U5258 ( .I(n3925), .ZN(n3446) );
  AOI22D0BWP U5259 ( .A1(op1[9]), .A2(n4672), .B1(op2[1]), .B2(n4671), .ZN(
        n3447) );
  NR2D0BWP U5260 ( .A1(n5759), .A2(n5758), .ZN(n3448) );
  MUX2ND0BWP U5261 ( .I0(n4845), .I1(n4844), .S(n4843), .ZN(n3449) );
  AOI22D0BWP U5262 ( .A1(n4689), .A2(n3448), .B1(n4690), .B2(n3449), .ZN(n3450) );
  OAI211D0BWP U5263 ( .A1(n3445), .A2(n3446), .B(n3447), .C(n3450), .ZN(
        result[9]) );
  AOI21D0BWP U5264 ( .A1(n4907), .A2(n4908), .B(n4871), .ZN(n3451) );
  NR2D0BWP U5265 ( .A1(n4955), .A2(n3451), .ZN(n4933) );
  CKND0BWP U5266 ( .I(n4548), .ZN(n3452) );
  MOAI22D0BWP U5267 ( .A1(n5416), .A2(n3452), .B1(n4549), .B2(n5414), .ZN(
        n3453) );
  AOI31D0BWP U5268 ( .A1(n3667), .A2(n5418), .A3(n5417), .B(n3453), .ZN(n3454)
         );
  IOA21D0BWP U5269 ( .A1(n3669), .A2(vectorToLoad[64]), .B(n3454), .ZN(N4281)
         );
  MUX2ND0BWP U5270 ( .I0(n3806), .I1(n3805), .S(nextInstrAddr[1]), .ZN(n3455)
         );
  MOAI22D0BWP U5271 ( .A1(n4643), .A2(n3939), .B1(n3455), .B2(n4061), .ZN(
        N4154) );
  AN2D0BWP U5272 ( .A1(\DP_OP_493J11_130_7648/n15 ), .A2(
        \DP_OP_493J11_130_7648/n44 ), .Z(\DP_OP_493J11_130_7648/n14 ) );
  INR2D0BWP U5273 ( .A1(n3773), .B1(\alu/N328 ), .ZN(n3864) );
  AN2D0BWP U5274 ( .A1(\DP_OP_493J11_130_7648/n18 ), .A2(
        \DP_OP_493J11_130_7648/n47 ), .Z(\DP_OP_493J11_130_7648/n17 ) );
  AN2D0BWP U5275 ( .A1(\DP_OP_493J11_130_7648/n22 ), .A2(
        \DP_OP_493J11_130_7648/n51 ), .Z(\DP_OP_493J11_130_7648/n21 ) );
  AN2D0BWP U5276 ( .A1(\DP_OP_493J11_130_7648/n26 ), .A2(
        \DP_OP_493J11_130_7648/n55 ), .Z(\DP_OP_493J11_130_7648/n25 ) );
  MUX2ND0BWP U5277 ( .I0(n4702), .I1(n4704), .S(n4237), .ZN(n3456) );
  CKND2D0BWP U5278 ( .A1(\intadd_34/SUM[1] ), .A2(n3456), .ZN(n4275) );
  AN2D0BWP U5279 ( .A1(\DP_OP_487J11_125_9213/n25 ), .A2(
        \DP_OP_487J11_125_9213/n54 ), .Z(\DP_OP_487J11_125_9213/n24 ) );
  AN2D0BWP U5280 ( .A1(\DP_OP_487J11_125_9213/n20 ), .A2(
        \DP_OP_487J11_125_9213/n49 ), .Z(\DP_OP_487J11_125_9213/n19 ) );
  INR2D0BWP U5281 ( .A1(N1470), .B1(n4351), .ZN(n4142) );
  INR2D0BWP U5282 ( .A1(n4146), .B1(n4097), .ZN(n4637) );
  MOAI22D0BWP U5283 ( .A1(n4803), .A2(n4801), .B1(n4800), .B2(n4799), .ZN(
        \mult_x_153/n140 ) );
  MOAI22D0BWP U5284 ( .A1(n4793), .A2(n4791), .B1(n5555), .B2(n4790), .ZN(
        \mult_x_153/n129 ) );
  CKND0BWP U5285 ( .I(n5709), .ZN(n3457) );
  AOI32D0BWP U5286 ( .A1(n5710), .A2(n5714), .A3(n3457), .B1(n5713), .B2(n5714), .ZN(n5728) );
  OAI21D0BWP U5287 ( .A1(n4464), .A2(n4463), .B(n3897), .ZN(n3458) );
  AOI211D0BWP U5288 ( .A1(n4464), .A2(n4463), .B(n5784), .C(n3458), .ZN(n3459)
         );
  AOI22D0BWP U5289 ( .A1(\alu/N684 ), .A2(n4657), .B1(n4659), .B2(n3459), .ZN(
        n3460) );
  AN3D0BWP U5290 ( .A1(n4460), .A2(n5704), .A3(n3460), .Z(n4656) );
  CKND0BWP U5291 ( .I(n4471), .ZN(n3461) );
  OA211D1BWP U5292 ( .A1(n4698), .A2(n5296), .B(n5295), .C(n3461), .Z(n4534)
         );
  CKND2D0BWP U5293 ( .A1(n4919), .A2(n4632), .ZN(n3462) );
  NR4D0BWP U5294 ( .A1(n4915), .A2(n4953), .A3(n4387), .A4(n3462), .ZN(n3463)
         );
  CKND0BWP U5295 ( .I(n4888), .ZN(n3464) );
  CKND0BWP U5296 ( .I(n4890), .ZN(n3465) );
  AOI221D0BWP U5297 ( .A1(n4890), .A2(n3464), .B1(n3465), .B2(n4888), .C(n4389), .ZN(n3466) );
  ND4D0BWP U5298 ( .A1(n4889), .A2(n4385), .A3(n4386), .A4(n3466), .ZN(n3467)
         );
  OAI31D0BWP U5299 ( .A1(n4633), .A2(n4891), .A3(n3467), .B(n4390), .ZN(n3468)
         );
  NR3D0BWP U5300 ( .A1(n4962), .A2(n3463), .A3(n3468), .ZN(n4967) );
  AOI22D0BWP U5301 ( .A1(n5233), .A2(vectorData2[180]), .B1(n5231), .B2(
        vectorData2[116]), .ZN(n3469) );
  AOI22D0BWP U5302 ( .A1(n5230), .A2(vectorData2[164]), .B1(n3601), .B2(
        vectorData2[36]), .ZN(n3470) );
  AOI22D0BWP U5303 ( .A1(n5232), .A2(vectorData2[148]), .B1(n5229), .B2(
        vectorData2[244]), .ZN(n3471) );
  CKND2D0BWP U5304 ( .A1(n3470), .A2(n3471), .ZN(n3472) );
  AOI21D0BWP U5305 ( .A1(vectorData2[196]), .A2(n5227), .B(n3472), .ZN(n3473)
         );
  AOI22D0BWP U5306 ( .A1(n5228), .A2(vectorData2[212]), .B1(n5226), .B2(
        vectorData2[132]), .ZN(n3474) );
  AOI31D0BWP U5307 ( .A1(n3469), .A2(n3473), .A3(n3474), .B(n3661), .ZN(n3475)
         );
  AOI22D0BWP U5308 ( .A1(n4694), .A2(vectorData2[228]), .B1(n4683), .B2(
        vectorData2[100]), .ZN(n3476) );
  AOI22D0BWP U5309 ( .A1(n4685), .A2(vectorData2[20]), .B1(n4684), .B2(
        vectorData2[84]), .ZN(n3477) );
  AOI22D0BWP U5310 ( .A1(n4681), .A2(vectorData2[4]), .B1(n4682), .B2(
        vectorData2[68]), .ZN(n3478) );
  AOI22D0BWP U5311 ( .A1(n4688), .A2(scalarData2[4]), .B1(n4686), .B2(
        vectorData2[52]), .ZN(n3479) );
  ND4D0BWP U5312 ( .A1(n3476), .A2(n3477), .A3(n3478), .A4(n3479), .ZN(n3480)
         );
  AO211D0BWP U5313 ( .A1(n3928), .A2(instrIn[4]), .B(n3475), .C(n3480), .Z(
        N4196) );
  NR2D0BWP U5314 ( .A1(n4989), .A2(nextInstrAddr[15]), .ZN(n3481) );
  AOI21D0BWP U5315 ( .A1(nextInstrAddr[14]), .A2(n4641), .B(n4391), .ZN(n3482)
         );
  AOI21D0BWP U5316 ( .A1(n4641), .A2(n3481), .B(n3482), .ZN(n3483) );
  OAI211D0BWP U5317 ( .A1(n3939), .A2(n6037), .B(n5998), .C(n3483), .ZN(N4169)
         );
  INR2D0BWP U5318 ( .A1(n3766), .B1(\alu/N337 ), .ZN(n3772) );
  AN2D0BWP U5319 ( .A1(\DP_OP_493J11_130_7648/n14 ), .A2(
        \DP_OP_493J11_130_7648/n43 ), .Z(\DP_OP_493J11_130_7648/n13 ) );
  AN2D0BWP U5320 ( .A1(\DP_OP_493J11_130_7648/n19 ), .A2(
        \DP_OP_493J11_130_7648/n48 ), .Z(\DP_OP_493J11_130_7648/n18 ) );
  AN2D0BWP U5321 ( .A1(\DP_OP_493J11_130_7648/n23 ), .A2(
        \DP_OP_493J11_130_7648/n52 ), .Z(\DP_OP_493J11_130_7648/n22 ) );
  INR2D0BWP U5322 ( .A1(\DP_OP_493J11_130_7648/n56 ), .B1(n5793), .ZN(
        \DP_OP_493J11_130_7648/n26 ) );
  AN2D0BWP U5323 ( .A1(\DP_OP_487J11_125_9213/n16 ), .A2(
        \DP_OP_487J11_125_9213/n45 ), .Z(\DP_OP_487J11_125_9213/n15 ) );
  AN2D0BWP U5324 ( .A1(\DP_OP_487J11_125_9213/n22 ), .A2(
        \DP_OP_487J11_125_9213/n51 ), .Z(\DP_OP_487J11_125_9213/n21 ) );
  AN2D0BWP U5325 ( .A1(\DP_OP_487J11_125_9213/n26 ), .A2(
        \DP_OP_487J11_125_9213/n55 ), .Z(\DP_OP_487J11_125_9213/n25 ) );
  AN2D0BWP U5326 ( .A1(\DP_OP_487J11_125_9213/n19 ), .A2(
        \DP_OP_487J11_125_9213/n48 ), .Z(\DP_OP_487J11_125_9213/n18 ) );
  AOI21D0BWP U5327 ( .A1(N1473), .A2(n4091), .B(N1475), .ZN(n3484) );
  CKND0BWP U5328 ( .I(N1477), .ZN(n3485) );
  OAI32D0BWP U5329 ( .A1(N1478), .A2(N1476), .A3(n3484), .B1(n3485), .B2(N1478), .ZN(n3486) );
  IAO21D0BWP U5330 ( .A1(N1479), .A2(n3486), .B(N1480), .ZN(n4101) );
  MOAI22D0BWP U5331 ( .A1(n4789), .A2(n5554), .B1(n4796), .B2(n4788), .ZN(
        \mult_x_153/n127 ) );
  INR2D0BWP U5332 ( .A1(n4463), .B1(n5711), .ZN(n4465) );
  IND3D0BWP U5333 ( .A1(func[2]), .B1(n1), .B2(n3487), .ZN(n3740) );
  CKND0BWP U5334 ( .I(func[3]), .ZN(n3487) );
  INR2D0BWP U5335 ( .A1(n4090), .B1(n4089), .ZN(n4146) );
  INR3D0BWP U5336 ( .A1(n3787), .B1(n3663), .B2(state[3]), .ZN(n3720) );
  AO21D0BWP U5337 ( .A1(n4673), .A2(n5747), .B(n5732), .Z(n3488) );
  AOI32D0BWP U5338 ( .A1(n5733), .A2(n5758), .A3(n3488), .B1(n5731), .B2(n5758), .ZN(n5745) );
  AOI32D0BWP U5339 ( .A1(n3871), .A2(n3869), .A3(n4410), .B1(n3870), .B2(n3869), .ZN(n3489) );
  OAI21D0BWP U5340 ( .A1(n4411), .A2(\intadd_35/SUM[1] ), .B(n3489), .ZN(n5777) );
  IND2D0BWP U5341 ( .A1(n6040), .B1(n5997), .ZN(N4211) );
  ND4D0BWP U5342 ( .A1(n8058), .A2(n8057), .A3(n8056), .A4(n8055), .ZN(n3490)
         );
  AOI22D0BWP U5343 ( .A1(n5233), .A2(vectorData1[190]), .B1(n5187), .B2(n3490), 
        .ZN(n3491) );
  AOI22D0BWP U5344 ( .A1(n5230), .A2(vectorData1[174]), .B1(n5186), .B2(
        vectorData1[78]), .ZN(n3492) );
  ND4D0BWP U5345 ( .A1(n7994), .A2(n7993), .A3(n7992), .A4(n7991), .ZN(n3493)
         );
  ND4D0BWP U5346 ( .A1(n5112), .A2(n5113), .A3(n5114), .A4(n5115), .ZN(n3494)
         );
  AOI21D0BWP U5347 ( .A1(n5228), .A2(n3493), .B(n3494), .ZN(n3495) );
  AOI22D0BWP U5348 ( .A1(n5232), .A2(vectorData1[158]), .B1(n5185), .B2(
        vectorData1[94]), .ZN(n3496) );
  AN4D0BWP U5349 ( .A1(n3491), .A2(n3492), .A3(n3495), .A4(n3496), .Z(n3497)
         );
  AOI22D0BWP U5350 ( .A1(n8278), .A2(\srf/regTable[0][14] ), .B1(n8280), .B2(
        \srf/regTable[2][14] ), .ZN(n3498) );
  AOI22D0BWP U5351 ( .A1(n8284), .A2(\srf/regTable[3][14] ), .B1(n8282), .B2(
        \srf/regTable[1][14] ), .ZN(n3499) );
  AOI22D0BWP U5352 ( .A1(n8285), .A2(\srf/regTable[4][14] ), .B1(n8286), .B2(
        \srf/regTable[6][14] ), .ZN(n3500) );
  AOI22D0BWP U5353 ( .A1(n8288), .A2(\srf/regTable[7][14] ), .B1(n8287), .B2(
        \srf/regTable[5][14] ), .ZN(n3501) );
  ND4D0BWP U5354 ( .A1(n3498), .A2(n3499), .A3(n3500), .A4(n3501), .ZN(n3502)
         );
  AOI22D0BWP U5355 ( .A1(n3581), .A2(\vrf/regTable[0][14] ), .B1(n3572), .B2(
        \vrf/regTable[2][14] ), .ZN(n3503) );
  AOI22D0BWP U5356 ( .A1(n3579), .A2(\vrf/regTable[1][14] ), .B1(n3575), .B2(
        \vrf/regTable[3][14] ), .ZN(n3504) );
  AOI22D0BWP U5357 ( .A1(n3574), .A2(\vrf/regTable[4][14] ), .B1(n3570), .B2(
        \vrf/regTable[6][14] ), .ZN(n3505) );
  AOI22D0BWP U5358 ( .A1(n3576), .A2(\vrf/regTable[5][14] ), .B1(n3567), .B2(
        \vrf/regTable[7][14] ), .ZN(n3506) );
  ND4D0BWP U5359 ( .A1(n3503), .A2(n3504), .A3(n3505), .A4(n3506), .ZN(n3507)
         );
  AOI22D0BWP U5360 ( .A1(n4073), .A2(n3502), .B1(n4072), .B2(n3507), .ZN(n3508) );
  CKND2D0BWP U5361 ( .A1(n4071), .A2(Addr[14]), .ZN(n3509) );
  OAI211D0BWP U5362 ( .A1(n4070), .A2(n3497), .B(n3508), .C(n3509), .ZN(N4190)
         );
  AOI22D0BWP U5363 ( .A1(n5231), .A2(vectorData2[123]), .B1(n5227), .B2(
        vectorData2[203]), .ZN(n3510) );
  AOI22D0BWP U5364 ( .A1(n5230), .A2(vectorData2[171]), .B1(n5229), .B2(
        vectorData2[251]), .ZN(n3511) );
  AOI22D0BWP U5365 ( .A1(n5226), .A2(vectorData2[139]), .B1(n5233), .B2(
        vectorData2[187]), .ZN(n3512) );
  AOI22D0BWP U5366 ( .A1(n5232), .A2(vectorData2[155]), .B1(n5228), .B2(
        vectorData2[219]), .ZN(n3513) );
  AN4D0BWP U5367 ( .A1(n3510), .A2(n3511), .A3(n3512), .A4(n3513), .Z(n3514)
         );
  AOI22D0BWP U5368 ( .A1(n4688), .A2(scalarData2[11]), .B1(n4681), .B2(
        vectorData2[11]), .ZN(n3515) );
  AOI22D0BWP U5369 ( .A1(n4682), .A2(vectorData2[75]), .B1(n4685), .B2(
        vectorData2[27]), .ZN(n3516) );
  AOI22D0BWP U5370 ( .A1(n4684), .A2(vectorData2[91]), .B1(n4686), .B2(
        vectorData2[59]), .ZN(n3517) );
  AOI22D0BWP U5371 ( .A1(n4687), .A2(vectorData2[43]), .B1(n4683), .B2(
        vectorData2[107]), .ZN(n3518) );
  ND4D0BWP U5372 ( .A1(n3515), .A2(n3516), .A3(n3517), .A4(n3518), .ZN(n3519)
         );
  AOI21D0BWP U5373 ( .A1(n4694), .A2(vectorData2[235]), .B(n3519), .ZN(n3520)
         );
  OAI211D0BWP U5374 ( .A1(n3661), .A2(n3514), .B(n3792), .C(n3520), .ZN(N4203)
         );
  CKND0BWP U5375 ( .I(vectorToLoad[192]), .ZN(n3521) );
  CKND0BWP U5376 ( .I(n5416), .ZN(n3522) );
  AOI22D0BWP U5377 ( .A1(n5415), .A2(n5414), .B1(n4534), .B2(n3522), .ZN(n3523) );
  OAI211D0BWP U5378 ( .A1(n3670), .A2(n3521), .B(n3523), .C(n4535), .ZN(n3524)
         );
  AO31D0BWP U5379 ( .A1(n4625), .A2(n5418), .A3(n5417), .B(n3524), .Z(N4410)
         );
  CKND0BWP U5380 ( .I(n4991), .ZN(n3525) );
  CKND0BWP U5381 ( .I(cycles[4]), .ZN(n3526) );
  AOI221D0BWP U5382 ( .A1(n4991), .A2(cycles[4]), .B1(n3525), .B2(n3526), .C(
        n4574), .ZN(N4175) );
  INR3D0BWP U5383 ( .A1(n4641), .B1(nextInstrAddr[14]), .B2(n4064), .ZN(n3527)
         );
  AOI211D0BWP U5384 ( .A1(result[14]), .A2(n4066), .B(n3527), .C(n4065), .ZN(
        n3528) );
  OAI21D0BWP U5385 ( .A1(n4641), .A2(n4989), .B(n3528), .ZN(N4168) );
  AN2D0BWP U5386 ( .A1(\DP_OP_493J11_130_7648/n17 ), .A2(
        \DP_OP_493J11_130_7648/n46 ), .Z(\DP_OP_493J11_130_7648/n16 ) );
  AN2D0BWP U5387 ( .A1(\DP_OP_493J11_130_7648/n21 ), .A2(
        \DP_OP_493J11_130_7648/n50 ), .Z(\DP_OP_493J11_130_7648/n20 ) );
  AN2D0BWP U5388 ( .A1(\DP_OP_493J11_130_7648/n25 ), .A2(
        \DP_OP_493J11_130_7648/n54 ), .Z(\DP_OP_493J11_130_7648/n24 ) );
  INR2D0BWP U5389 ( .A1(n3865), .B1(n3866), .ZN(\intadd_35/B[1] ) );
  INR2D0BWP U5390 ( .A1(n4182), .B1(\intadd_34/SUM[1] ), .ZN(n4274) );
  AN2D0BWP U5391 ( .A1(\DP_OP_487J11_125_9213/n56 ), .A2(\C1/Z_0 ), .Z(
        \DP_OP_487J11_125_9213/n26 ) );
  AN2D0BWP U5392 ( .A1(\DP_OP_487J11_125_9213/n24 ), .A2(
        \DP_OP_487J11_125_9213/n53 ), .Z(\DP_OP_487J11_125_9213/n23 ) );
  AN2D0BWP U5393 ( .A1(\DP_OP_487J11_125_9213/n21 ), .A2(
        \DP_OP_487J11_125_9213/n50 ), .Z(\DP_OP_487J11_125_9213/n20 ) );
  AN2D0BWP U5394 ( .A1(\DP_OP_487J11_125_9213/n18 ), .A2(
        \DP_OP_487J11_125_9213/n47 ), .Z(\DP_OP_487J11_125_9213/n17 ) );
  AN2D0BWP U5395 ( .A1(\DP_OP_487J11_125_9213/n15 ), .A2(
        \DP_OP_487J11_125_9213/n44 ), .Z(\DP_OP_487J11_125_9213/n14 ) );
  CKND0BWP U5396 ( .I(N1472), .ZN(n3529) );
  OAI21D0BWP U5397 ( .A1(n4093), .A2(n3529), .B(n4094), .ZN(n3530) );
  AOI21D0BWP U5398 ( .A1(n4096), .A2(n3530), .B(n4095), .ZN(n4143) );
  IND2D0BWP U5399 ( .A1(n4055), .B1(n4056), .ZN(n5793) );
  CKND0BWP U5400 ( .I(n4462), .ZN(n3531) );
  AOI21D0BWP U5401 ( .A1(n4460), .A2(n3531), .B(n4461), .ZN(n3532) );
  CKND2D0BWP U5402 ( .A1(n4674), .A2(n4458), .ZN(n3533) );
  CKND2D0BWP U5403 ( .A1(n4459), .A2(n3533), .ZN(n3534) );
  OAI211D0BWP U5404 ( .A1(n4459), .A2(n3533), .B(n5739), .C(n3534), .ZN(n3535)
         );
  OAI21D0BWP U5405 ( .A1(n5739), .A2(n3532), .B(n3535), .ZN(n5738) );
  IND2D0BWP U5406 ( .A1(n3727), .B1(n3728), .ZN(n3712) );
  AOI22D0BWP U5407 ( .A1(n5802), .A2(\intadd_33/SUM[3] ), .B1(n5801), .B2(
        \intadd_33/SUM[2] ), .ZN(n3536) );
  CKND0BWP U5408 ( .I(n3925), .ZN(n3537) );
  AOI22D0BWP U5409 ( .A1(op2[3]), .A2(n4672), .B1(op1[3]), .B2(n4671), .ZN(
        n3538) );
  NR2D0BWP U5410 ( .A1(n5754), .A2(n5727), .ZN(n3539) );
  MUX2ND0BWP U5411 ( .I0(n4856), .I1(n5556), .S(n4855), .ZN(n3540) );
  AOI22D0BWP U5412 ( .A1(n4689), .A2(n3539), .B1(n4690), .B2(n3540), .ZN(n3541) );
  OAI211D0BWP U5413 ( .A1(n3536), .A2(n3537), .B(n3538), .C(n3541), .ZN(
        result[3]) );
  CKND0BWP U5414 ( .I(n4896), .ZN(n3542) );
  CKND0BWP U5415 ( .I(n4903), .ZN(n3543) );
  AOI32D0BWP U5416 ( .A1(n4634), .A2(n3542), .A3(n3543), .B1(n4896), .B2(n4156), .ZN(n4911) );
  OAI31D0BWP U5417 ( .A1(n4633), .A2(n4964), .A3(n4965), .B(n4963), .ZN(n3544)
         );
  AOI32D0BWP U5418 ( .A1(n4966), .A2(n4639), .A3(n4632), .B1(n3544), .B2(n4639), .ZN(n3545) );
  AOI32D0BWP U5419 ( .A1(\intadd_34/A[3] ), .A2(n3545), .A3(n4474), .B1(n4967), 
        .B2(n3545), .ZN(N1824) );
  AOI22D0BWP U5420 ( .A1(n5227), .A2(vectorData2[206]), .B1(n5232), .B2(
        vectorData2[158]), .ZN(n3546) );
  AOI22D0BWP U5421 ( .A1(n5233), .A2(vectorData2[190]), .B1(n5226), .B2(
        vectorData2[142]), .ZN(n3547) );
  AOI22D0BWP U5422 ( .A1(n5230), .A2(vectorData2[174]), .B1(n5228), .B2(
        vectorData2[222]), .ZN(n3548) );
  AOI22D0BWP U5423 ( .A1(n5229), .A2(vectorData2[254]), .B1(n5231), .B2(
        vectorData2[126]), .ZN(n3549) );
  AN4D0BWP U5424 ( .A1(n3546), .A2(n3547), .A3(n3548), .A4(n3549), .Z(n3550)
         );
  AOI22D0BWP U5425 ( .A1(n4688), .A2(scalarData2[14]), .B1(n4685), .B2(
        vectorData2[30]), .ZN(n3551) );
  AOI22D0BWP U5426 ( .A1(n4682), .A2(vectorData2[78]), .B1(n4694), .B2(
        vectorData2[238]), .ZN(n3552) );
  AOI22D0BWP U5427 ( .A1(n4684), .A2(vectorData2[94]), .B1(n4683), .B2(
        vectorData2[110]), .ZN(n3553) );
  AOI22D0BWP U5428 ( .A1(n4686), .A2(vectorData2[62]), .B1(n4687), .B2(
        vectorData2[46]), .ZN(n3554) );
  ND4D0BWP U5429 ( .A1(n3551), .A2(n3552), .A3(n3553), .A4(n3554), .ZN(n3555)
         );
  AOI21D0BWP U5430 ( .A1(n4681), .A2(vectorData2[14]), .B(n3555), .ZN(n3556)
         );
  OAI211D0BWP U5431 ( .A1(n3661), .A2(n3550), .B(n3792), .C(n3556), .ZN(N4206)
         );
  OR2D0BWP U5432 ( .A1(WR), .A2(RD), .Z(N4133) );
  CKND2D0BWP U5433 ( .A1(cycles[2]), .A2(n4992), .ZN(n3557) );
  AOI211D0BWP U5434 ( .A1(n3675), .A2(n3557), .B(n4991), .C(n4574), .ZN(N4174)
         );
  INR2D0BWP U5435 ( .A1(n3932), .B1(n3861), .ZN(n3558) );
  OAI211D0BWP U5436 ( .A1(nextInstrAddr[12]), .A2(n3558), .B(n4061), .C(n4062), 
        .ZN(n3559) );
  OAI211D0BWP U5437 ( .A1(n3939), .A2(\intadd_34/A[1] ), .B(n5998), .C(n3559), 
        .ZN(N4166) );
  NR2D3BWP U5438 ( .A1(n3663), .A2(state[3]), .ZN(n3719) );
  ND2D1BWP U5439 ( .A1(n3562), .A2(n3707), .ZN(n3560) );
  CKND2BWP U5440 ( .I(n3560), .ZN(n4068) );
  ND3D3BWP U5441 ( .A1(n156), .A2(n3712), .A3(n4616), .ZN(n3713) );
  CKND12BWP U5442 ( .I(Reset), .ZN(n156) );
  CKBD4BWP U5443 ( .I(n7115), .Z(n3574) );
  CKBD4BWP U5444 ( .I(n7108), .Z(n3581) );
  CKBD4BWP U5445 ( .I(n6080), .Z(n3577) );
  CKBD4BWP U5446 ( .I(n6073), .Z(n3580) );
  INVD1BWP U5447 ( .I(n5793), .ZN(n4612) );
  IND2D2BWP U5448 ( .A1(n3611), .B1(n3605), .ZN(n3613) );
  ND2D4BWP U5449 ( .A1(n3563), .A2(n3664), .ZN(n3783) );
  CKND2BWP U5450 ( .I(n3564), .ZN(n3565) );
  NR3D0BWP U5451 ( .A1(n3793), .A2(Reset), .A3(n4393), .ZN(n4066) );
  ND2D8BWP U5452 ( .A1(n6039), .A2(n4623), .ZN(n6063) );
  CKND3BWP U5453 ( .I(n4505), .ZN(n4535) );
  IND2D1BWP U5454 ( .A1(state[3]), .B1(n3562), .ZN(n3611) );
  OAI21D1BWP U5455 ( .A1(n3721), .A2(n3783), .B(n3609), .ZN(n3722) );
  CKBD1BWP U5456 ( .I(\intadd_34/n1 ), .Z(\intadd_34/CO ) );
  INVD1BWP U5457 ( .I(\intadd_34/SUM[1] ), .ZN(n4254) );
  CKND1BWP U5458 ( .I(\intadd_34/SUM[0] ), .ZN(n4237) );
  INR2D1BWP U5459 ( .A1(n3613), .B1(n3722), .ZN(n3602) );
  INR2D2BWP U5460 ( .A1(n3565), .B1(n3606), .ZN(n3605) );
  NR2XD0BWP U5461 ( .A1(n6074), .A2(\vrf/N14 ), .ZN(n6075) );
  BUFFD6BWP U5462 ( .I(n6082), .Z(n3569) );
  BUFFD6BWP U5463 ( .I(n6077), .Z(n3571) );
  ND3D1BWP U5464 ( .A1(n3663), .A2(n4573), .A3(state[3]), .ZN(n3608) );
  NR2D1BWP U5465 ( .A1(n3732), .A2(n4573), .ZN(n3717) );
  AOI21D1BWP U5466 ( .A1(n3702), .A2(n3701), .B(n3783), .ZN(n3703) );
  BUFFD6BWP U5467 ( .I(n7117), .Z(n3576) );
  CKND0BWP U5468 ( .I(n4573), .ZN(n3598) );
  NR3D1BWP U5469 ( .A1(\vrf/N12 ), .A2(\vrf/N13 ), .A3(n4622), .ZN(n8210) );
  NR3D1BWP U5470 ( .A1(\vrf/N9 ), .A2(\vrf/N10 ), .A3(n4619), .ZN(n8285) );
  BUFFD6BWP U5471 ( .I(n7112), .Z(n3579) );
  NR2XD0BWP U5472 ( .A1(n6078), .A2(\vrf/N14 ), .ZN(n6079) );
  CKND2D1BWP U5473 ( .A1(n3726), .A2(n3718), .ZN(n3702) );
  NR3D1BWP U5474 ( .A1(\vrf/N14 ), .A2(\vrf/N12 ), .A3(\vrf/N13 ), .ZN(n8203)
         );
  NR3D1BWP U5475 ( .A1(\vrf/N11 ), .A2(\vrf/N9 ), .A3(\vrf/N10 ), .ZN(n8278)
         );
  CKND2D1BWP U5476 ( .A1(n3726), .A2(n3700), .ZN(n3701) );
  NR2D0BWP U5477 ( .A1(n4558), .A2(code[0]), .ZN(n4623) );
  INVD1BWP U5478 ( .I(n3746), .ZN(n4561) );
  NR2D2BWP U5479 ( .A1(n5509), .A2(n5817), .ZN(n5415) );
  BUFFD1BWP U5480 ( .I(n4628), .Z(n3667) );
  NR2D1BWP U5481 ( .A1(n5509), .A2(cycles[3]), .ZN(n4505) );
  CKND1BWP U5482 ( .I(op1[9]), .ZN(n3680) );
  CKBD2BWP U5483 ( .I(n4630), .Z(n3582) );
  CKND2D0BWP U5484 ( .A1(code[2]), .A2(n3698), .ZN(n3786) );
  CKND1BWP U5485 ( .I(code[1]), .ZN(n4697) );
  INVD0BWP U5486 ( .I(code[0]), .ZN(n3699) );
  AN2XD1BWP U5487 ( .A1(n4548), .A2(n4547), .Z(n3649) );
  CKND2D1BWP U5488 ( .A1(n4398), .A2(n4471), .ZN(N4215) );
  NR2D0BWP U5489 ( .A1(n4394), .A2(n3782), .ZN(RD) );
  NR2D0BWP U5490 ( .A1(n4393), .A2(n3562), .ZN(n4395) );
  ND2D1BWP U5491 ( .A1(n3562), .A2(n3681), .ZN(n3697) );
  NR2D1BWP U5492 ( .A1(n3679), .A2(n5417), .ZN(n4992) );
  NR2D2BWP U5493 ( .A1(state[1]), .A2(state[3]), .ZN(n3681) );
  INVD1BWP U5494 ( .I(state[3]), .ZN(n3726) );
  INVD1BWP U5495 ( .I(cycles[0]), .ZN(n3679) );
  INVD1BWP U5496 ( .I(cycles[4]), .ZN(n4698) );
  CKND1BWP U5497 ( .I(cycles[1]), .ZN(n5417) );
  INVD1BWP U5498 ( .I(cycles[2]), .ZN(n5812) );
  MAOI22D0BWP U5499 ( .A1(n4125), .A2(n4124), .B1(n4123), .B2(n4122), .ZN(
        n4131) );
  MAOI22D0BWP U5500 ( .A1(N1483), .A2(n4360), .B1(n4887), .B2(n4358), .ZN(
        n4356) );
  AN4D1BWP U5501 ( .A1(n4115), .A2(n4114), .A3(n4113), .A4(n4112), .Z(n4116)
         );
  MAOI22D0BWP U5502 ( .A1(N1478), .A2(n4351), .B1(N1481), .B2(n4107), .ZN(
        n4346) );
  CKXOR2D1BWP U5503 ( .A1(\DP_OP_487J11_125_9213/n1 ), .A2(\C1/Z_0 ), .Z(N1483) );
  CKXOR2D0BWP U5504 ( .A1(\DP_OP_487J11_125_9213/n14 ), .A2(
        \DP_OP_487J11_125_9213/n43 ), .Z(N1470) );
  MAOI22D0BWP U5505 ( .A1(n4694), .A2(vectorData2[224]), .B1(n5129), .B2(n3661), .ZN(n3756) );
  MAOI22D0BWP U5506 ( .A1(n4694), .A2(vectorData2[227]), .B1(n5156), .B2(n3661), .ZN(n3820) );
  AN4D1BWP U5507 ( .A1(n5155), .A2(n5154), .A3(n5153), .A4(n5152), .Z(n5156)
         );
  AN4D1BWP U5508 ( .A1(n5128), .A2(n5127), .A3(n5126), .A4(n5125), .Z(n5129)
         );
  AN3D1BWP U5509 ( .A1(nextInstrAddr[9]), .A2(n3929), .A3(nextInstrAddr[10]), 
        .Z(n3932) );
  AN3D1BWP U5510 ( .A1(nextInstrAddr[8]), .A2(nextInstrAddr[7]), .A3(n3922), 
        .Z(n3929) );
  AN3D1BWP U5511 ( .A1(n3858), .A2(nextInstrAddr[5]), .A3(nextInstrAddr[6]), 
        .Z(n3922) );
  AN3D1BWP U5512 ( .A1(n3838), .A2(nextInstrAddr[3]), .A3(nextInstrAddr[4]), 
        .Z(n3858) );
  AN3D1BWP U5513 ( .A1(n3805), .A2(nextInstrAddr[1]), .A3(nextInstrAddr[2]), 
        .Z(n3838) );
  OAI31D1BWP U5514 ( .A1(\srf/N15 ), .A2(n138), .A3(n8202), .B(n156), .ZN(
        \srf/N53 ) );
  OAI31D1BWP U5515 ( .A1(\srf/N15 ), .A2(n3651), .A3(n8202), .B(n156), .ZN(
        \srf/N55 ) );
  OAI31D1BWP U5516 ( .A1(n138), .A2(n3637), .A3(n8202), .B(n156), .ZN(
        \srf/N36 ) );
  OAI31D1BWP U5517 ( .A1(n3637), .A2(n3651), .A3(n8202), .B(n156), .ZN(
        \srf/N54 ) );
  OAI31D1BWP U5518 ( .A1(\srf/N15 ), .A2(n138), .A3(\srf/N17 ), .B(n156), .ZN(
        \srf/N57 ) );
  OAI31D1BWP U5519 ( .A1(\srf/N15 ), .A2(\srf/N17 ), .A3(n3651), .B(n156), 
        .ZN(\srf/N59 ) );
  OAI31D1BWP U5520 ( .A1(\srf/N17 ), .A2(n3637), .A3(n3651), .B(n156), .ZN(
        \srf/N58 ) );
  OAI31D1BWP U5521 ( .A1(n138), .A2(\srf/N17 ), .A3(n3637), .B(n156), .ZN(
        \srf/N56 ) );
  IND2D1BWP U5522 ( .A1(n6001), .B1(n6000), .ZN(n6038) );
  MAOI22D0BWP U5523 ( .A1(n4320), .A2(n4326), .B1(n4324), .B2(n4260), .ZN(
        n4207) );
  OR4XD1BWP U5524 ( .A1(n4696), .A2(n5247), .A3(Reset), .A4(n4060), .Z(N4162)
         );
  OA222D1BWP U5525 ( .A1(n4237), .A2(n4702), .B1(n4254), .B2(n4182), .C1(n4234), .C2(n4704), .Z(n4300) );
  MAOI22D0BWP U5526 ( .A1(n4228), .A2(result[0]), .B1(n4705), .B2(n4237), .ZN(
        n4249) );
  MAOI22D0BWP U5527 ( .A1(n4227), .A2(n4169), .B1(\intadd_34/SUM[0] ), .B2(
        n4708), .ZN(n4225) );
  AO31D1BWP U5528 ( .A1(n4689), .A2(n4656), .A3(n5753), .B(n3902), .Z(
        result[7]) );
  CKND1BWP U5529 ( .I(result[1]), .ZN(n4643) );
  AN4D1BWP U5530 ( .A1(n3777), .A2(n3776), .A3(n3775), .A4(n3774), .Z(n3778)
         );
  CKXOR2D1BWP U5531 ( .A1(\DP_OP_493J11_130_7648/n1 ), .A2(n4612), .Z(
        \alu/N339 ) );
  CKXOR2D0BWP U5532 ( .A1(\DP_OP_493J11_130_7648/n14 ), .A2(
        \DP_OP_493J11_130_7648/n43 ), .Z(\alu/N326 ) );
  XNR2D1BWP U5533 ( .A1(result[15]), .A2(n4336), .ZN(\C1/Z_0 ) );
  AOI31D0BWP U5534 ( .A1(n4642), .A2(n4542), .A3(n4474), .B(n4541), .ZN(n4545)
         );
  MAOI22D0BWP U5535 ( .A1(n4002), .A2(n4035), .B1(n4006), .B2(n4033), .ZN(
        n3996) );
  INR3D0BWP U5536 ( .A1(n3613), .B1(n3704), .B2(n3703), .ZN(n3705) );
  MAOI22D0BWP U5537 ( .A1(n4002), .A2(n4032), .B1(n4006), .B2(n4031), .ZN(
        n3997) );
  MAOI22D0BWP U5538 ( .A1(n4048), .A2(n4035), .B1(n4034), .B2(n4033), .ZN(
        n4036) );
  MAOI22D0BWP U5539 ( .A1(n4048), .A2(n4032), .B1(n4034), .B2(n4031), .ZN(
        n4037) );
  NR2D1BWP U5540 ( .A1(n3696), .A2(n3695), .ZN(n3706) );
  MAOI22D0BWP U5541 ( .A1(n4731), .A2(n4751), .B1(n4751), .B2(n4730), .ZN(
        n4734) );
  MAOI22D0BWP U5542 ( .A1(n4649), .A2(n4740), .B1(n4741), .B2(n4649), .ZN(
        n4755) );
  MAOI22D0BWP U5543 ( .A1(n4750), .A2(n4751), .B1(n3959), .B2(n3960), .ZN(
        n3983) );
  MAOI22D0BWP U5544 ( .A1(n4649), .A2(n4721), .B1(n4720), .B2(n4649), .ZN(
        n4733) );
  MAOI22D0BWP U5545 ( .A1(n4730), .A2(n4751), .B1(n3961), .B2(n3960), .ZN(
        n3982) );
  MAOI22D0BWP U5546 ( .A1(n4752), .A2(n4751), .B1(n4751), .B2(n4750), .ZN(
        n4756) );
  MAOI22D0BWP U5547 ( .A1(n3652), .A2(n4726), .B1(n4725), .B2(n3652), .ZN(
        n4731) );
  MAOI22D0BWP U5548 ( .A1(n3652), .A2(n4746), .B1(n4745), .B2(n3652), .ZN(
        n4752) );
  BUFFD3BWP U5549 ( .I(n7110), .Z(n3594) );
  BUFFD3BWP U5550 ( .I(n7118), .Z(n3595) );
  NR2D1BWP U5551 ( .A1(Reset), .A2(n4573), .ZN(n3710) );
  BUFFD3BWP U5552 ( .I(n7116), .Z(n3596) );
  MAOI22D0BWP U5553 ( .A1(n5555), .A2(n4795), .B1(n4774), .B2(n4793), .ZN(
        n4776) );
  BUFFD3BWP U5554 ( .I(n7114), .Z(n3599) );
  MAOI22D0BWP U5555 ( .A1(n5563), .A2(n5572), .B1(n5567), .B2(n5562), .ZN(
        n5586) );
  INR2D1BWP U5556 ( .A1(n4623), .B1(n4468), .ZN(n6040) );
  CKND1BWP U5557 ( .I(n4558), .ZN(n4554) );
  OA21D1BWP U5558 ( .A1(op2[10]), .A2(op1[10]), .B(n3950), .Z(n5622) );
  CKND2D0BWP U5559 ( .A1(code[0]), .A2(n3712), .ZN(n4553) );
  OAI21D1BWP U5560 ( .A1(n5561), .A2(n4666), .B(n5613), .ZN(n4820) );
  OAI21D1BWP U5561 ( .A1(n4832), .A2(n4662), .B(n5614), .ZN(n4808) );
  NR2XD0BWP U5562 ( .A1(n4568), .A2(n4566), .ZN(n4570) );
  IND2D1BWP U5563 ( .A1(n3610), .B1(n3720), .ZN(n3609) );
  CKND2D1BWP U5564 ( .A1(n3698), .A2(n4561), .ZN(n4558) );
  OAI21D1BWP U5565 ( .A1(n4478), .A2(n4695), .B(n4552), .ZN(n4070) );
  CKND0BWP U5566 ( .I(n3728), .ZN(n3689) );
  CKMUX2D1BWP U5567 ( .I0(n5811), .I1(n4552), .S(n137), .Z(n3692) );
  AOI211D0BWP U5568 ( .A1(code[0]), .A2(n4992), .B(cycles[4]), .C(n3728), .ZN(
        n3687) );
  CKND1BWP U5569 ( .I(n3666), .ZN(n3665) );
  CKND1BWP U5570 ( .I(op1[3]), .ZN(n5561) );
  CKND1BWP U5571 ( .I(op1[5]), .ZN(n4832) );
  AOI21D1BWP U5572 ( .A1(n3786), .A2(n4567), .B(n3788), .ZN(n4073) );
  NR2XD0BWP U5573 ( .A1(n4568), .A2(n4567), .ZN(n4569) );
  CKND1BWP U5574 ( .I(n4551), .ZN(n4552) );
  INVD2BWP U5575 ( .I(n4631), .ZN(n3670) );
  CKND1BWP U5576 ( .I(op1[7]), .ZN(n5605) );
  INR3D0BWP U5577 ( .A1(func[2]), .B1(func[3]), .B2(n3739), .ZN(n4672) );
  NR3D0BWP U5578 ( .A1(func[3]), .A2(n3734), .A3(n3738), .ZN(n4671) );
  NR2XD0BWP U5579 ( .A1(n3740), .A2(func[0]), .ZN(n4689) );
  NR2D0BWP U5580 ( .A1(n4697), .A2(n3786), .ZN(n3746) );
  AN4D1BWP U5581 ( .A1(n3740), .A2(n3739), .A3(n3738), .A4(n3737), .Z(n4690)
         );
  NR3D0BWP U5582 ( .A1(func[3]), .A2(func[2]), .A3(n3739), .ZN(n4691) );
  CKBD2BWP U5583 ( .I(n4630), .Z(n3600) );
  INR2D1BWP U5584 ( .A1(n5249), .B1(n4397), .ZN(n4631) );
  NR2XD0BWP U5585 ( .A1(n4473), .A2(n5812), .ZN(n4628) );
  NR3D0BWP U5586 ( .A1(n132), .A2(n5812), .A3(n4543), .ZN(n4625) );
  CKND0BWP U5587 ( .I(N4215), .ZN(n4397) );
  CKND1BWP U5588 ( .I(code[3]), .ZN(n3698) );
  CKND0BWP U5589 ( .I(code[2]), .ZN(n3684) );
  AN2XD1BWP U5590 ( .A1(n4548), .A2(n4470), .Z(n3650) );
  ND2D1BWP U5591 ( .A1(n4534), .A2(n3617), .ZN(n4405) );
  CKND1BWP U5592 ( .I(n4477), .ZN(n4538) );
  INR3D0BWP U5593 ( .A1(n4698), .B1(n5296), .B2(n4398), .ZN(n4408) );
  NR2XD0BWP U5594 ( .A1(n3784), .A2(Reset), .ZN(n4061) );
  NR2XD0BWP U5595 ( .A1(n4468), .A2(Reset), .ZN(n6039) );
  AN4D1BWP U5596 ( .A1(n5830), .A2(n4564), .A3(n4563), .A4(n4562), .Z(n4565)
         );
  NR2XD2BWP U5597 ( .A1(n3783), .A2(n3711), .ZN(n4616) );
  CKND1BWP U5598 ( .I(n3682), .ZN(n4542) );
  ND2D1BWP U5599 ( .A1(RD), .A2(n3562), .ZN(n4471) );
  CKND2D0BWP U5600 ( .A1(n4395), .A2(n4394), .ZN(n4468) );
  NR2XD1BWP U5601 ( .A1(n4996), .A2(n4998), .ZN(n5227) );
  NR2XD1BWP U5602 ( .A1(n4995), .A2(n4993), .ZN(n5231) );
  NR2XD1BWP U5603 ( .A1(n4997), .A2(n4994), .ZN(n5228) );
  CKND1BWP U5604 ( .I(n4992), .ZN(n5811) );
  NR2XD1BWP U5605 ( .A1(n4995), .A2(n4998), .ZN(n5233) );
  AOI21D0BWP U5606 ( .A1(n3679), .A2(n5417), .B(n4992), .ZN(n5292) );
  INVD1BWP U5607 ( .I(n3616), .ZN(n3601) );
  NR2XD1BWP U5608 ( .A1(n4999), .A2(n4998), .ZN(n5230) );
  NR2XD1BWP U5609 ( .A1(n4997), .A2(n4998), .ZN(n5232) );
  NR2XD1BWP U5610 ( .A1(n4995), .A2(n4994), .ZN(n5229) );
  INVD1BWP U5611 ( .I(n3681), .ZN(n3782) );
  INR2XD0BWP U5612 ( .A1(n3663), .B1(n3612), .ZN(n3707) );
  NR2D1BWP U5613 ( .A1(n3726), .A2(state[1]), .ZN(n3716) );
  IND2D0BWP U5614 ( .A1(n3612), .B1(state[1]), .ZN(n4393) );
  CKND2D0BWP U5615 ( .A1(cycles[0]), .A2(n5287), .ZN(n5290) );
  CKND2D0BWP U5616 ( .A1(n5807), .A2(n5251), .ZN(n5249) );
  NR2D0BWP U5617 ( .A1(n5251), .A2(n5293), .ZN(n5291) );
  CKND0BWP U5618 ( .I(n5813), .ZN(n5293) );
  CKND2D0BWP U5619 ( .A1(n137), .A2(n5818), .ZN(n5282) );
  NR2D0BWP U5620 ( .A1(cycles[4]), .A2(cycles[3]), .ZN(n5807) );
  NR3D0BWP U5621 ( .A1(cycles[2]), .A2(cycles[0]), .A3(cycles[1]), .ZN(n5251)
         );
  NR2XD0BWP U5622 ( .A1(cycles[2]), .A2(cycles[1]), .ZN(n5294) );
  CKND0BWP U5623 ( .I(cycles[3]), .ZN(n3675) );
  NR3D1BWP U5624 ( .A1(\srf/N17 ), .A2(\srf/N15 ), .A3(n3651), .ZN(n8127) );
  NR3D1BWP U5625 ( .A1(\srf/N15 ), .A2(n3651), .A3(n8202), .ZN(n8134) );
  AOI21D1BWP U5626 ( .A1(n3602), .A2(n3603), .B(Reset), .ZN(N153) );
  AOI21D1BWP U5627 ( .A1(n3725), .A2(n3604), .B(n3660), .ZN(n3603) );
  IND2D1BWP U5628 ( .A1(n3607), .B1(n3694), .ZN(n3695) );
  INVD1BWP U5629 ( .I(n3719), .ZN(n3711) );
  ND2D1BWP U5630 ( .A1(n3719), .A2(n3718), .ZN(n3721) );
  ND3D1BWP U5631 ( .A1(n3719), .A2(n3787), .A3(n156), .ZN(n3708) );
  NR3D2BWP U5632 ( .A1(n3697), .A2(n3664), .A3(n4573), .ZN(n3704) );
  INVD1BWP U5633 ( .I(n4068), .ZN(n3614) );
  CKND2BWP U5634 ( .I(n3670), .ZN(n3669) );
  CKND2BWP U5635 ( .I(n3670), .ZN(n3668) );
  MAOI22D0BWP U5636 ( .A1(n4477), .A2(DataIn[0]), .B1(n5299), .B2(n4473), .ZN(
        n4476) );
  CKND2D0BWP U5637 ( .A1(n6039), .A2(n5999), .ZN(n6001) );
  ND2D1BWP U5638 ( .A1(code[0]), .A2(n4392), .ZN(n6000) );
  MAOI222D1BWP U5639 ( .A(n5581), .B(n5580), .C(n5579), .ZN(n5582) );
  CKND2BWP U5640 ( .I(n5692), .ZN(n4650) );
  NR2XD1BWP U5641 ( .A1(n4993), .A2(n4996), .ZN(n5226) );
  ND2D1BWP U5642 ( .A1(code[0]), .A2(n3727), .ZN(n4567) );
  NR3D1BWP U5643 ( .A1(n5818), .A2(n5817), .A3(n5816), .ZN(n5982) );
  NR3D1BWP U5644 ( .A1(n5818), .A2(n5817), .A3(n5815), .ZN(n5983) );
  CKND6BWP U5645 ( .I(n3664), .ZN(n4394) );
  CKND4BWP U5646 ( .I(n3564), .ZN(n3664) );
  MOAI22D0BWP U5647 ( .A1(n5513), .A2(n3666), .B1(n4534), .B2(n5512), .ZN(
        n4479) );
  MOAI22D0BWP U5648 ( .A1(n5538), .A2(n3666), .B1(n4534), .B2(n5537), .ZN(
        n4504) );
  ND2D1BWP U5649 ( .A1(n4571), .A2(n156), .ZN(N4209) );
  INVD1BWP U5650 ( .I(n4571), .ZN(N4208) );
  INVD1BWP U5651 ( .I(n5511), .ZN(n5513) );
  INVD1BWP U5652 ( .I(n5410), .ZN(n5506) );
  INVD1BWP U5653 ( .I(n5412), .ZN(n5510) );
  ND2D1BWP U5654 ( .A1(n4933), .A2(n4967), .ZN(n4909) );
  INVD1BWP U5655 ( .I(vectorToLoad[245]), .ZN(n4515) );
  INVD1BWP U5656 ( .I(vectorToLoad[246]), .ZN(n4517) );
  INVD1BWP U5657 ( .I(vectorToLoad[247]), .ZN(n4519) );
  INVD1BWP U5658 ( .I(vectorToLoad[248]), .ZN(n4521) );
  INVD1BWP U5659 ( .I(vectorToLoad[249]), .ZN(n4523) );
  AN2XD1BWP U5660 ( .A1(n5294), .A2(n5403), .Z(n3630) );
  INVD1BWP U5661 ( .I(vectorToLoad[250]), .ZN(n4525) );
  AN2XD1BWP U5662 ( .A1(n5294), .A2(n5357), .Z(n3623) );
  INVD1BWP U5663 ( .I(vectorToLoad[251]), .ZN(n4527) );
  AN2XD1BWP U5664 ( .A1(n5294), .A2(n5406), .Z(n3631) );
  INVD1BWP U5665 ( .I(vectorToLoad[252]), .ZN(n4529) );
  AN2XD1BWP U5666 ( .A1(n5294), .A2(n5408), .Z(n3632) );
  INVD1BWP U5667 ( .I(vectorToLoad[253]), .ZN(n4531) );
  AN2XD1BWP U5668 ( .A1(n5294), .A2(n5410), .Z(n3633) );
  INVD1BWP U5669 ( .I(vectorToLoad[254]), .ZN(n4533) );
  INVD1BWP U5670 ( .I(vectorToLoad[255]), .ZN(n4537) );
  AN2XD1BWP U5671 ( .A1(n5294), .A2(n5400), .Z(n3629) );
  INVD1BWP U5672 ( .I(vectorToLoad[244]), .ZN(n4513) );
  ND2D1BWP U5673 ( .A1(n4066), .A2(result[2]), .ZN(n3815) );
  ND2D1BWP U5674 ( .A1(n4066), .A2(result[5]), .ZN(n3848) );
  ND2D1BWP U5675 ( .A1(n4066), .A2(result[7]), .ZN(n3907) );
  ND2D1BWP U5676 ( .A1(n4066), .A2(result[13]), .ZN(n3935) );
  ND2D1BWP U5677 ( .A1(n5462), .A2(n4549), .ZN(n4544) );
  INVD1BWP U5678 ( .I(vectorToLoad[16]), .ZN(n4546) );
  INVD1BWP U5679 ( .I(n4066), .ZN(n3939) );
  ND2D1BWP U5680 ( .A1(n4066), .A2(result[11]), .ZN(n3933) );
  AN2XD1BWP U5681 ( .A1(n5294), .A2(n5352), .Z(n3622) );
  ND2D1BWP U5682 ( .A1(n4066), .A2(result[9]), .ZN(n3930) );
  ND2D1BWP U5683 ( .A1(n3562), .A2(n3664), .ZN(n3793) );
  AN2XD1BWP U5684 ( .A1(n5294), .A2(n5341), .Z(n3621) );
  ND2D1BWP U5685 ( .A1(n4534), .A2(n5514), .ZN(n4409) );
  INVD1BWP U5686 ( .I(vectorToLoad[228]), .ZN(n4481) );
  AN2XD1BWP U5687 ( .A1(n5294), .A2(n5394), .Z(n3626) );
  INVD1BWP U5688 ( .I(vectorToLoad[229]), .ZN(n4483) );
  INVD1BWP U5689 ( .I(vectorToLoad[230]), .ZN(n4485) );
  INVD1BWP U5690 ( .I(vectorToLoad[231]), .ZN(n4487) );
  INVD1BWP U5691 ( .I(vectorToLoad[232]), .ZN(n4489) );
  INVD1BWP U5692 ( .I(vectorToLoad[233]), .ZN(n4491) );
  INVD1BWP U5693 ( .I(vectorToLoad[234]), .ZN(n4493) );
  INVD1BWP U5694 ( .I(vectorToLoad[235]), .ZN(n4495) );
  AN2XD1BWP U5695 ( .A1(n5294), .A2(n5396), .Z(n3627) );
  INVD1BWP U5696 ( .I(vectorToLoad[236]), .ZN(n4497) );
  INVD1BWP U5697 ( .I(vectorToLoad[237]), .ZN(n4499) );
  AN2XD1BWP U5698 ( .A1(n5293), .A2(n5328), .Z(n3648) );
  INVD1BWP U5699 ( .I(vectorToLoad[238]), .ZN(n4501) );
  AN2XD1BWP U5700 ( .A1(n5293), .A2(n5330), .Z(n3636) );
  INVD1BWP U5701 ( .I(vectorToLoad[239]), .ZN(n4503) );
  INVD1BWP U5702 ( .I(n4540), .ZN(n4629) );
  ND2D1BWP U5703 ( .A1(n4548), .A2(n3617), .ZN(n4540) );
  INVD1BWP U5704 ( .I(n5536), .ZN(n5538) );
  AN2XD1BWP U5705 ( .A1(n5294), .A2(n5412), .Z(n3634) );
  AN2XD1BWP U5706 ( .A1(n5294), .A2(n5387), .Z(n3620) );
  INVD1BWP U5707 ( .I(vectorToLoad[241]), .ZN(n4507) );
  AN2XD1BWP U5708 ( .A1(n5294), .A2(n5398), .Z(n3628) );
  AN2XD1BWP U5709 ( .A1(n5294), .A2(n5389), .Z(n3624) );
  INVD1BWP U5710 ( .I(vectorToLoad[242]), .ZN(n4509) );
  ND2D1BWP U5711 ( .A1(n4956), .A2(n4967), .ZN(n4906) );
  AN2XD1BWP U5712 ( .A1(n5294), .A2(n5391), .Z(n3625) );
  INVD1BWP U5713 ( .I(n4625), .ZN(n3666) );
  INVD1BWP U5714 ( .I(vectorToLoad[243]), .ZN(n4511) );
  ND2D1BWP U5715 ( .A1(n4688), .A2(scalarData2[10]), .ZN(n3796) );
  INVD1BWP U5716 ( .I(n3944), .ZN(n3797) );
  AN2XD1BWP U5717 ( .A1(n4548), .A2(n5514), .Z(n3654) );
  INVD1BWP U5718 ( .I(vectorData2[114]), .ZN(n5143) );
  ND2D1BWP U5719 ( .A1(n4404), .A2(n4406), .ZN(N4346) );
  ND2D1BWP U5720 ( .A1(n5299), .A2(cycles[3]), .ZN(n4402) );
  INVD1BWP U5721 ( .I(nextInstrAddr[0]), .ZN(n3806) );
  INVD1BWP U5722 ( .I(vectorData2[129]), .ZN(n5132) );
  AN2XD1BWP U5723 ( .A1(n5293), .A2(n5308), .Z(n3635) );
  AN2XD1BWP U5724 ( .A1(n5293), .A2(n5310), .Z(n3639) );
  INVD1BWP U5725 ( .I(nextInstrAddr[11]), .ZN(n3861) );
  ND2D1BWP U5726 ( .A1(n5297), .A2(n5287), .ZN(n5416) );
  INVD1BWP U5727 ( .I(n5370), .ZN(n5297) );
  INVD1BWP U5728 ( .I(nextInstrAddr[13]), .ZN(n4063) );
  INVD1BWP U5729 ( .I(n4061), .ZN(n4064) );
  ND2D1BWP U5730 ( .A1(n4061), .A2(nextInstrAddr[14]), .ZN(n4989) );
  INVD1BWP U5731 ( .I(n4983), .ZN(n4067) );
  ND2D1BWP U5732 ( .A1(n4061), .A2(nextInstrAddr[15]), .ZN(n4391) );
  ND2D1BWP U5733 ( .A1(n4980), .A2(n4981), .ZN(n4983) );
  INVD1BWP U5734 ( .I(n4978), .ZN(n4981) );
  INVD1BWP U5735 ( .I(n4975), .ZN(n4976) );
  ND2D1BWP U5736 ( .A1(result[9]), .A2(n4974), .ZN(n4975) );
  ND2D1BWP U5737 ( .A1(n3903), .A2(result[7]), .ZN(n3918) );
  ND2D1BWP U5738 ( .A1(n4973), .A2(result[5]), .ZN(n3854) );
  ND2D1BWP U5739 ( .A1(cycles[4]), .A2(n4970), .ZN(n4972) );
  INVD1BWP U5740 ( .I(n5231), .ZN(n3674) );
  INVD1BWP U5741 ( .I(vectorData2[124]), .ZN(n5203) );
  INVD1BWP U5742 ( .I(n5240), .ZN(n3792) );
  INVD1BWP U5743 ( .I(n5419), .ZN(n4470) );
  ND2D1BWP U5744 ( .A1(n137), .A2(n5287), .ZN(n5288) );
  INVD1BWP U5745 ( .I(n5314), .ZN(n5437) );
  INVD1BWP U5746 ( .I(n5316), .ZN(n5440) );
  AN2XD1BWP U5747 ( .A1(n5293), .A2(n5320), .Z(n3644) );
  INVD1BWP U5748 ( .I(n5318), .ZN(n5443) );
  INVD1BWP U5749 ( .I(n5320), .ZN(n5446) );
  INVD1BWP U5750 ( .I(n5322), .ZN(n5449) );
  INVD1BWP U5751 ( .I(n5324), .ZN(n5452) );
  INVD1BWP U5752 ( .I(n5326), .ZN(n5455) );
  AN2XD1BWP U5753 ( .A1(n5293), .A2(n5322), .Z(n3645) );
  INVD1BWP U5754 ( .I(n5328), .ZN(n5458) );
  INVD1BWP U5755 ( .I(n5387), .ZN(n5467) );
  INVD1BWP U5756 ( .I(n5389), .ZN(n5470) );
  AN2XD1BWP U5757 ( .A1(n5293), .A2(n5324), .Z(n3646) );
  INVD1BWP U5758 ( .I(n5391), .ZN(n5473) );
  INVD1BWP U5759 ( .I(n5394), .ZN(n5479) );
  INVD1BWP U5760 ( .I(n5396), .ZN(n5482) );
  INVD1BWP U5761 ( .I(n5398), .ZN(n5485) );
  INVD1BWP U5762 ( .I(n5400), .ZN(n5488) );
  AN2XD1BWP U5763 ( .A1(n5293), .A2(n5326), .Z(n3647) );
  INVD1BWP U5764 ( .I(n5403), .ZN(n5494) );
  INVD1BWP U5765 ( .I(n5406), .ZN(n5500) );
  INVD1BWP U5766 ( .I(n5312), .ZN(n5434) );
  INVD1BWP U5767 ( .I(n5330), .ZN(n5461) );
  ND2D1BWP U5768 ( .A1(result[1]), .A2(n4399), .ZN(n5335) );
  AN2XD1BWP U5769 ( .A1(n5293), .A2(n5312), .Z(n3640) );
  ND2D1BWP U5770 ( .A1(result[2]), .A2(n4399), .ZN(n5337) );
  ND2D1BWP U5771 ( .A1(result[3]), .A2(n4399), .ZN(n5339) );
  INVD1BWP U5772 ( .I(n5341), .ZN(n5476) );
  ND2D1BWP U5773 ( .A1(result[5]), .A2(n4399), .ZN(n5344) );
  ND2D1BWP U5774 ( .A1(result[6]), .A2(n4399), .ZN(n5346) );
  ND2D1BWP U5775 ( .A1(result[7]), .A2(n4399), .ZN(n5348) );
  ND2D1BWP U5776 ( .A1(n4073), .A2(scalarData1[4]), .ZN(n3831) );
  ND2D1BWP U5777 ( .A1(n5186), .A2(vectorData1[68]), .ZN(n3827) );
  ND2D1BWP U5778 ( .A1(n5041), .A2(n5043), .ZN(n3829) );
  ND2D1BWP U5779 ( .A1(n3601), .A2(vectorData1[36]), .ZN(n5043) );
  AN2XD1BWP U5780 ( .A1(n5293), .A2(n5314), .Z(n3641) );
  ND2D1BWP U5781 ( .A1(result[8]), .A2(n4399), .ZN(n5350) );
  INVD1BWP U5782 ( .I(Addr[3]), .ZN(n3823) );
  INVD1BWP U5783 ( .I(n5352), .ZN(n5491) );
  INVD1BWP U5784 ( .I(n5464), .ZN(n5289) );
  ND2D1BWP U5785 ( .A1(DataIn[0]), .A2(n3679), .ZN(n5464) );
  ND2D1BWP U5786 ( .A1(result[10]), .A2(n4399), .ZN(n5355) );
  INVD1BWP U5787 ( .I(Addr[2]), .ZN(n3808) );
  INVD1BWP U5788 ( .I(n5357), .ZN(n5497) );
  ND2D1BWP U5789 ( .A1(result[12]), .A2(n4399), .ZN(n5360) );
  AN2XD1BWP U5790 ( .A1(n5293), .A2(n5316), .Z(n3642) );
  ND2D1BWP U5791 ( .A1(result[13]), .A2(n4399), .ZN(n5362) );
  ND2D1BWP U5792 ( .A1(result[14]), .A2(n4399), .ZN(n5364) );
  INVD1BWP U5793 ( .I(Addr[0]), .ZN(n3789) );
  ND2D1BWP U5794 ( .A1(n4627), .A2(n3675), .ZN(n4406) );
  INVD1BWP U5795 ( .I(n4405), .ZN(n4626) );
  NR2XD0BWP U5796 ( .A1(n5812), .A2(cycles[1]), .ZN(n5287) );
  ND2D1BWP U5797 ( .A1(result[15]), .A2(n4399), .ZN(n5366) );
  ND2D1BWP U5798 ( .A1(cycles[0]), .A2(n5254), .ZN(n5334) );
  INVD1BWP U5799 ( .I(n4642), .ZN(n5286) );
  ND2D1BWP U5800 ( .A1(DataIn[0]), .A2(cycles[0]), .ZN(n5370) );
  INVD1BWP U5801 ( .I(n5301), .ZN(n5517) );
  INVD1BWP U5802 ( .I(n5304), .ZN(n5520) );
  AN2XD1BWP U5803 ( .A1(n5293), .A2(n5318), .Z(n3643) );
  INVD1BWP U5804 ( .I(n5306), .ZN(n5523) );
  INVD1BWP U5805 ( .I(n4408), .ZN(n4543) );
  INVD1BWP U5806 ( .I(n5308), .ZN(n5428) );
  INVD1BWP U5807 ( .I(n5310), .ZN(n5431) );
  INVD1BWP U5808 ( .I(n5292), .ZN(n4990) );
  INVD1BWP U5809 ( .I(n5408), .ZN(n5503) );
  ND2D1BWP U5810 ( .A1(n3911), .A2(n3910), .ZN(N4200) );
  ND2D1BWP U5811 ( .A1(n4681), .A2(vectorData2[5]), .ZN(n3842) );
  INVD1BWP U5812 ( .I(n3928), .ZN(n3844) );
  ND2D1BWP U5813 ( .A1(n3883), .A2(n3747), .ZN(n3928) );
  ND2D1BWP U5814 ( .A1(n3946), .A2(n3945), .ZN(N4201) );
  INVD1BWP U5815 ( .I(vectorData2[143]), .ZN(n5236) );
  ND2D1BWP U5816 ( .A1(n5418), .A2(n5254), .ZN(n5299) );
  AN2XD1BWP U5817 ( .A1(n137), .A2(result[0]), .Z(n5418) );
  INVD1BWP U5818 ( .I(DataIn[12]), .ZN(n5279) );
  INVD1BWP U5819 ( .I(DataIn[13]), .ZN(n5280) );
  INVD1BWP U5820 ( .I(DataIn[15]), .ZN(n5283) );
  ND2D1BWP U5821 ( .A1(n4478), .A2(n5250), .ZN(n4539) );
  ND2D1BWP U5822 ( .A1(n137), .A2(n5254), .ZN(n5302) );
  INVD1BWP U5823 ( .I(n132), .ZN(n5298) );
  INVD1BWP U5824 ( .I(n5249), .ZN(n4474) );
  INVD1BWP U5825 ( .I(n4572), .ZN(n4466) );
  INVD1BWP U5826 ( .I(n3830), .ZN(n4071) );
  ND2D1BWP U5827 ( .A1(n4616), .A2(n3787), .ZN(n3830) );
  NR3D1BWP U5828 ( .A1(\vrf/N9 ), .A2(\vrf/N10 ), .A3(n4619), .ZN(n7115) );
  ND2D1BWP U5829 ( .A1(\vrf/N9 ), .A2(\vrf/N10 ), .ZN(n7113) );
  ND2D1BWP U5830 ( .A1(\vrf/N9 ), .A2(n4617), .ZN(n7111) );
  ND2D1BWP U5831 ( .A1(\vrf/N10 ), .A2(n4618), .ZN(n7109) );
  NR3D1BWP U5832 ( .A1(\vrf/N11 ), .A2(\vrf/N9 ), .A3(\vrf/N10 ), .ZN(n7108)
         );
  INVD1BWP U5833 ( .I(\vrf/N11 ), .ZN(n4619) );
  ND2D1BWP U5834 ( .A1(\vrf/N9 ), .A2(\vrf/N10 ), .ZN(n8283) );
  ND2D1BWP U5835 ( .A1(\vrf/N9 ), .A2(n4617), .ZN(n8281) );
  INVD1BWP U5836 ( .I(\vrf/N10 ), .ZN(n4617) );
  ND2D1BWP U5837 ( .A1(\vrf/N10 ), .A2(n4618), .ZN(n8279) );
  INVD1BWP U5838 ( .I(\vrf/N9 ), .ZN(n4618) );
  INVD1BWP U5839 ( .I(instrIn[6]), .ZN(n4556) );
  INVD1BWP U5840 ( .I(n4616), .ZN(n3788) );
  INVD1BWP U5841 ( .I(n4953), .ZN(n4954) );
  ND2D1BWP U5842 ( .A1(n4957), .A2(n4949), .ZN(n4947) );
  ND2D1BWP U5843 ( .A1(n4700), .A2(n4942), .ZN(n4943) );
  INVD1BWP U5844 ( .I(n4933), .ZN(n4940) );
  ND2D1BWP U5845 ( .A1(n4932), .A2(n4931), .ZN(n4938) );
  ND2D1BWP U5846 ( .A1(n4941), .A2(n4935), .ZN(n4952) );
  INVD1BWP U5847 ( .I(n4911), .ZN(n4929) );
  ND2D1BWP U5848 ( .A1(n4156), .A2(n4155), .ZN(n4930) );
  INVD1BWP U5849 ( .I(n4914), .ZN(n4927) );
  INVD1BWP U5850 ( .I(n4757), .ZN(\mult_x_153/n41 ) );
  INVD1BWP U5851 ( .I(n4763), .ZN(\mult_x_153/n46 ) );
  INVD1BWP U5852 ( .I(n4773), .ZN(\mult_x_153/n87 ) );
  INVD1BWP U5853 ( .I(n4963), .ZN(n4924) );
  ND2D1BWP U5854 ( .A1(n4961), .A2(n4948), .ZN(n4963) );
  INVD1BWP U5855 ( .I(n4164), .ZN(n4165) );
  ND2D1BWP U5856 ( .A1(n4910), .A2(n4913), .ZN(n4936) );
  INVD1BWP U5857 ( .I(n4892), .ZN(n4161) );
  INVD1BWP U5858 ( .I(n4912), .ZN(n4910) );
  INVD1BWP U5859 ( .I(n4966), .ZN(n4961) );
  INVD1BWP U5860 ( .I(n4639), .ZN(n4962) );
  ND2D1BWP U5861 ( .A1(scalarToLoad[12]), .A2(scalarToLoad[11]), .ZN(n4076) );
  INVD1BWP U5862 ( .I(n4934), .ZN(n4387) );
  INVD1BWP U5863 ( .I(n4955), .ZN(n4965) );
  INVD1BWP U5864 ( .I(n4904), .ZN(n4869) );
  ND2D1BWP U5865 ( .A1(n4922), .A2(n4889), .ZN(n4964) );
  INVD1BWP U5866 ( .I(n4915), .ZN(n4700) );
  ND2D1BWP U5867 ( .A1(n4879), .A2(n4889), .ZN(n4882) );
  ND2D1BWP U5868 ( .A1(n4878), .A2(n4890), .ZN(n4880) );
  ND2D1BWP U5869 ( .A1(n4376), .A2(n4375), .ZN(n4377) );
  ND2D1BWP U5870 ( .A1(N1483), .A2(n4863), .ZN(n4118) );
  INVD1BWP U5871 ( .I(n4884), .ZN(n4375) );
  INVD1BWP U5872 ( .I(n4877), .ZN(n4119) );
  ND2D1BWP U5873 ( .A1(n4368), .A2(n4367), .ZN(n4877) );
  INVD1BWP U5874 ( .I(n4635), .ZN(n4367) );
  INVD1BWP U5875 ( .I(n4886), .ZN(n4383) );
  INVD1BWP U5876 ( .I(n4873), .ZN(n4901) );
  INVD1BWP U5877 ( .I(n4872), .ZN(n4902) );
  ND2D1BWP U5878 ( .A1(n4349), .A2(n4152), .ZN(n4104) );
  ND2D1BWP U5879 ( .A1(N1479), .A2(n4342), .ZN(n4098) );
  ND2D1BWP U5880 ( .A1(n4873), .A2(n4872), .ZN(n4870) );
  ND2D1BWP U5881 ( .A1(n4373), .A2(n4141), .ZN(n4130) );
  INVD1BWP U5882 ( .I(n4345), .ZN(n4125) );
  ND2D1BWP U5883 ( .A1(n4349), .A2(n4352), .ZN(n4109) );
  ND2D1BWP U5884 ( .A1(N1480), .A2(n4342), .ZN(n4343) );
  INVD1BWP U5885 ( .I(n4122), .ZN(n4342) );
  ND2D1BWP U5886 ( .A1(n4359), .A2(n4636), .ZN(n4345) );
  ND2D1BWP U5887 ( .A1(N1480), .A2(N1479), .ZN(n4107) );
  INVD1BWP U5888 ( .I(n4637), .ZN(n4100) );
  ND2D1BWP U5889 ( .A1(n4634), .A2(n4896), .ZN(n4898) );
  INVD1BWP U5890 ( .I(n4126), .ZN(n4128) );
  ND2D1BWP U5891 ( .A1(n4159), .A2(n4160), .ZN(n4894) );
  ND2D1BWP U5892 ( .A1(N1470), .A2(n4102), .ZN(n4103) );
  INVD1BWP U5893 ( .I(n4101), .ZN(n4102) );
  INVD1BWP U5894 ( .I(n4370), .ZN(n4384) );
  ND2D1BWP U5895 ( .A1(n4636), .A2(n4352), .ZN(n4122) );
  INVD1BWP U5896 ( .I(n4359), .ZN(n4352) );
  ND2D1BWP U5897 ( .A1(n4337), .A2(n4370), .ZN(n4341) );
  ND2D1BWP U5898 ( .A1(N1482), .A2(n4374), .ZN(n4370) );
  INVD1BWP U5899 ( .I(n4373), .ZN(n4148) );
  ND2D1BWP U5900 ( .A1(n4090), .A2(n4089), .ZN(n4866) );
  ND2D1BWP U5901 ( .A1(n4376), .A2(n4362), .ZN(n4363) );
  ND2D1BWP U5902 ( .A1(n4360), .A2(n4351), .ZN(n4358) );
  INVD1BWP U5903 ( .I(n4355), .ZN(n4351) );
  INVD1BWP U5904 ( .I(n4120), .ZN(n4362) );
  INVD1BWP U5905 ( .I(n4887), .ZN(n4366) );
  ND2D1BWP U5906 ( .A1(n4338), .A2(n4337), .ZN(n4887) );
  ND2D1BWP U5907 ( .A1(n4096), .A2(n4094), .ZN(n4089) );
  ND2D1BWP U5908 ( .A1(n4091), .A2(n4092), .ZN(n4093) );
  INVD1BWP U5909 ( .I(N1473), .ZN(n4092) );
  INVD1BWP U5910 ( .I(N1474), .ZN(n4091) );
  INVD1BWP U5911 ( .I(n4376), .ZN(n4338) );
  INVD1BWP U5912 ( .I(N1483), .ZN(n4374) );
  INVD1BWP U5913 ( .I(n4273), .ZN(n4262) );
  INVD1BWP U5914 ( .I(n4319), .ZN(n4259) );
  INVD1BWP U5915 ( .I(n4267), .ZN(n4268) );
  INVD1BWP U5916 ( .I(n4299), .ZN(n4266) );
  INVD1BWP U5917 ( .I(n4255), .ZN(n4233) );
  INVD1BWP U5918 ( .I(n4249), .ZN(n4313) );
  INVD1BWP U5919 ( .I(n4323), .ZN(n4315) );
  ND2D1BWP U5920 ( .A1(\intadd_34/SUM[0] ), .A2(n4261), .ZN(n4321) );
  INVD1BWP U5921 ( .I(n4709), .ZN(n4261) );
  INVD1BWP U5922 ( .I(n4333), .ZN(n4322) );
  ND2D1BWP U5923 ( .A1(\intadd_34/SUM[3] ), .A2(n4253), .ZN(n4323) );
  ND2D1BWP U5924 ( .A1(n4638), .A2(n4240), .ZN(n4232) );
  INVD1BWP U5925 ( .I(scalarToLoad[0]), .ZN(n4240) );
  INVD1BWP U5926 ( .I(n4225), .ZN(n4281) );
  INVD1BWP U5927 ( .I(n4260), .ZN(n4246) );
  INVD1BWP U5928 ( .I(n4223), .ZN(n4279) );
  INVD1BWP U5929 ( .I(n4222), .ZN(n4280) );
  ND2D1BWP U5930 ( .A1(n4221), .A2(n4220), .ZN(n4306) );
  INVD1BWP U5931 ( .I(scalarToLoad[1]), .ZN(n4162) );
  ND2D1BWP U5932 ( .A1(n4329), .A2(n4216), .ZN(n4217) );
  ND2D1BWP U5933 ( .A1(\intadd_34/SUM[1] ), .A2(n4213), .ZN(n4269) );
  ND2D1BWP U5934 ( .A1(n4212), .A2(n4211), .ZN(n4299) );
  INVD1BWP U5935 ( .I(n4331), .ZN(n4218) );
  INVD1BWP U5936 ( .I(n4301), .ZN(n4271) );
  INVD1BWP U5937 ( .I(n4703), .ZN(n4208) );
  INVD1BWP U5938 ( .I(n4215), .ZN(n4210) );
  INVD1BWP U5939 ( .I(scalarToLoad[2]), .ZN(n4158) );
  ND2D1BWP U5940 ( .A1(n4254), .A2(n4253), .ZN(n4215) );
  ND2D1BWP U5941 ( .A1(n4711), .A2(n4254), .ZN(n4197) );
  INVD1BWP U5942 ( .I(n4272), .ZN(n4320) );
  ND2D1BWP U5943 ( .A1(\intadd_34/SUM[2] ), .A2(n4195), .ZN(n4272) );
  INVD1BWP U5944 ( .I(scalarToLoad[3]), .ZN(n4157) );
  INVD1BWP U5945 ( .I(n4285), .ZN(n4192) );
  INVD1BWP U5946 ( .I(scalarToLoad[4]), .ZN(n4154) );
  ND2D1BWP U5947 ( .A1(n4227), .A2(scalarToLoad[6]), .ZN(n4185) );
  IOA22D1BWP U5948 ( .B1(n4664), .B2(\intadd_34/CO ), .A1(scalarToLoad[5]), 
        .A2(\intadd_34/CO ), .ZN(\C2/Z_20 ) );
  INVD1BWP U5949 ( .I(n4226), .ZN(n4241) );
  INVD1BWP U5950 ( .I(scalarToLoad[6]), .ZN(n4133) );
  INVD1BWP U5951 ( .I(n4234), .ZN(n4180) );
  ND2D1BWP U5952 ( .A1(n4237), .A2(n4254), .ZN(n4234) );
  INVD1BWP U5953 ( .I(n4707), .ZN(n4196) );
  ND2D1BWP U5954 ( .A1(n4178), .A2(n4177), .ZN(n4205) );
  INVD1BWP U5955 ( .I(n4288), .ZN(n4188) );
  INVD1BWP U5956 ( .I(n4286), .ZN(n4191) );
  INVD1BWP U5957 ( .I(n4228), .ZN(n4200) );
  INVD1BWP U5958 ( .I(n4227), .ZN(n4202) );
  INVD1BWP U5959 ( .I(scalarToLoad[7]), .ZN(n4187) );
  INVD1BWP U5960 ( .I(scalarToLoad[8]), .ZN(n4106) );
  ND2D1BWP U5961 ( .A1(\intadd_34/CO ), .A2(n4242), .ZN(n4175) );
  INVD1BWP U5962 ( .I(scalarToLoad[9]), .ZN(n4088) );
  ND2D1BWP U5963 ( .A1(n4242), .A2(n3676), .ZN(n4176) );
  ND2D1BWP U5964 ( .A1(result[10]), .A2(n4167), .ZN(n4168) );
  INVD1BWP U5965 ( .I(n4638), .ZN(n4706) );
  INVD1BWP U5966 ( .I(n4169), .ZN(n4087) );
  INVD1BWP U5967 ( .I(\intadd_34/CO ), .ZN(n3676) );
  ND2D1BWP U5968 ( .A1(n4219), .A2(n4169), .ZN(n4181) );
  ND2D1BWP U5969 ( .A1(\intadd_34/A[3] ), .A2(n4085), .ZN(n4169) );
  INVD1BWP U5970 ( .I(n4201), .ZN(n4219) );
  INVD1BWP U5971 ( .I(n4193), .ZN(n4166) );
  ND2D1BWP U5972 ( .A1(n4195), .A2(n4253), .ZN(n4260) );
  INVD1BWP U5973 ( .I(\intadd_34/SUM[2] ), .ZN(n4253) );
  INVD1BWP U5974 ( .I(\intadd_34/SUM[3] ), .ZN(n4195) );
  ND2D1BWP U5975 ( .A1(n4179), .A2(n4254), .ZN(n4258) );
  INVD1BWP U5976 ( .I(n4170), .ZN(n4167) );
  ND2D1BWP U5977 ( .A1(n4638), .A2(n4237), .ZN(n4201) );
  ND2D1BWP U5978 ( .A1(result[10]), .A2(n3615), .ZN(\intadd_34/CI ) );
  ND2D1BWP U5979 ( .A1(scalarToLoad[1]), .A2(n4469), .ZN(n6005) );
  ND2D1BWP U5980 ( .A1(scalarToLoad[0]), .A2(n4469), .ZN(n6002) );
  ND2D1BWP U5981 ( .A1(scalarToLoad[15]), .A2(n4469), .ZN(n6035) );
  ND2D1BWP U5982 ( .A1(scalarToLoad[14]), .A2(n4469), .ZN(n6032) );
  ND2D1BWP U5983 ( .A1(scalarToLoad[13]), .A2(n4469), .ZN(n6030) );
  ND2D1BWP U5984 ( .A1(scalarToLoad[12]), .A2(n4469), .ZN(n6028) );
  ND2D1BWP U5985 ( .A1(scalarToLoad[11]), .A2(n4469), .ZN(n6026) );
  INVD1BWP U5986 ( .I(result[11]), .ZN(\intadd_34/A[0] ) );
  ND2D1BWP U5987 ( .A1(scalarToLoad[10]), .A2(n4469), .ZN(n6024) );
  INVD1BWP U5988 ( .I(result[10]), .ZN(n4699) );
  ND2D1BWP U5989 ( .A1(scalarToLoad[9]), .A2(n4469), .ZN(n6022) );
  INVD1BWP U5990 ( .I(result[9]), .ZN(n4651) );
  ND2D1BWP U5991 ( .A1(scalarToLoad[8]), .A2(n4469), .ZN(n6020) );
  INVD1BWP U5992 ( .I(result[8]), .ZN(n4652) );
  ND2D1BWP U5993 ( .A1(scalarToLoad[7]), .A2(n4469), .ZN(n6018) );
  INVD1BWP U5994 ( .I(result[7]), .ZN(n4655) );
  ND2D1BWP U5995 ( .A1(scalarToLoad[6]), .A2(n4469), .ZN(n6016) );
  ND2D1BWP U5996 ( .A1(scalarToLoad[5]), .A2(n4469), .ZN(n6014) );
  INVD1BWP U5997 ( .I(result[5]), .ZN(n4664) );
  ND2D1BWP U5998 ( .A1(scalarToLoad[4]), .A2(n4469), .ZN(n6012) );
  ND2D1BWP U5999 ( .A1(scalarToLoad[3]), .A2(n4469), .ZN(n6009) );
  ND2D1BWP U6000 ( .A1(scalarToLoad[2]), .A2(n4469), .ZN(n6007) );
  INVD1BWP U6001 ( .I(\srf/N17 ), .ZN(n8202) );
  ND2D1BWP U6002 ( .A1(\srf/N15 ), .A2(n3651), .ZN(n8132) );
  ND2D1BWP U6003 ( .A1(\srf/N15 ), .A2(n138), .ZN(n8130) );
  ND2D1BWP U6004 ( .A1(n3651), .A2(n3637), .ZN(n8128) );
  INVD1BWP U6005 ( .I(n5998), .ZN(n4065) );
  ND2D1BWP U6006 ( .A1(n5247), .A2(n156), .ZN(n5998) );
  INVD1BWP U6007 ( .I(n5997), .ZN(n5999) );
  ND2D1BWP U6008 ( .A1(n4689), .A2(\alu/N665 ), .ZN(n3741) );
  INVD1BWP U6009 ( .I(n5784), .ZN(n5785) );
  ND2D1BWP U6010 ( .A1(n4690), .A2(\alu/N1018 ), .ZN(n3742) );
  ND2D1BWP U6011 ( .A1(\alu/N1003 ), .A2(n3925), .ZN(n3743) );
  INVD1BWP U6012 ( .I(result[13]), .ZN(\intadd_34/A[2] ) );
  ND2D1BWP U6013 ( .A1(n5775), .A2(n5777), .ZN(n5781) );
  INVD1BWP U6014 ( .I(result[12]), .ZN(\intadd_34/A[1] ) );
  INVD1BWP U6015 ( .I(n5788), .ZN(n5776) );
  INVD1BWP U6016 ( .I(n5769), .ZN(n5762) );
  ND2D1BWP U6017 ( .A1(n4465), .A2(n4464), .ZN(n5782) );
  ND2D1BWP U6018 ( .A1(n5804), .A2(n5803), .ZN(\alu/N832 ) );
  ND2D1BWP U6019 ( .A1(n5674), .A2(n5673), .ZN(n5679) );
  ND2D1BWP U6020 ( .A1(n5686), .A2(n5685), .ZN(n5687) );
  ND2D1BWP U6021 ( .A1(n3652), .A2(n5665), .ZN(n5626) );
  INVD1BWP U6022 ( .I(n5680), .ZN(n5667) );
  INVD1BWP U6023 ( .I(n5678), .ZN(n5666) );
  ND2D1BWP U6024 ( .A1(n5623), .A2(n5794), .ZN(n5678) );
  ND2D1BWP U6025 ( .A1(n5802), .A2(n5623), .ZN(n5680) );
  ND2D1BWP U6026 ( .A1(n5668), .A2(n5669), .ZN(n5676) );
  ND2D1BWP U6027 ( .A1(n5622), .A2(n5648), .ZN(n5656) );
  INVD1BWP U6028 ( .I(n5625), .ZN(n5648) );
  ND2D1BWP U6029 ( .A1(n5638), .A2(n5637), .ZN(n5639) );
  ND2D1BWP U6030 ( .A1(n5795), .A2(n5693), .ZN(n5634) );
  INVD1BWP U6031 ( .I(n5649), .ZN(\intadd_36/B[2] ) );
  INVD1BWP U6032 ( .I(n5645), .ZN(n5673) );
  INVD1BWP U6033 ( .I(n5665), .ZN(n5636) );
  INVD1BWP U6034 ( .I(n5647), .ZN(n5655) );
  INVD1BWP U6035 ( .I(result[15]), .ZN(n6037) );
  INVD1BWP U6036 ( .I(n4712), .ZN(n4835) );
  INVD1BWP U6037 ( .I(result[3]), .ZN(n6011) );
  INVD1BWP U6038 ( .I(result[0]), .ZN(n6004) );
  ND2D1BWP U6039 ( .A1(\alu/N990 ), .A2(n3925), .ZN(n3915) );
  ND2D1BWP U6040 ( .A1(n4656), .A2(n5756), .ZN(n5759) );
  ND2D1BWP U6041 ( .A1(\alu/N989 ), .A2(n3925), .ZN(n3899) );
  ND2D1BWP U6042 ( .A1(n4849), .A2(n4848), .ZN(n4847) );
  ND2D1BWP U6043 ( .A1(n5761), .A2(n5749), .ZN(n5790) );
  ND2D1BWP U6044 ( .A1(n5748), .A2(n5747), .ZN(n5749) );
  INVD1BWP U6045 ( .I(n5745), .ZN(n5774) );
  INVD1BWP U6046 ( .I(n5772), .ZN(n5752) );
  ND2D1BWP U6047 ( .A1(n5735), .A2(n5734), .ZN(n5737) );
  INVD1BWP U6048 ( .I(n4673), .ZN(n5748) );
  INVD1BWP U6049 ( .I(n5730), .ZN(n5758) );
  ND2D1BWP U6050 ( .A1(n5728), .A2(n5727), .ZN(n5732) );
  AN2XD1BWP U6051 ( .A1(n5736), .A2(n5740), .Z(n5733) );
  ND2D1BWP U6052 ( .A1(n5757), .A2(n5755), .ZN(n5731) );
  INVD1BWP U6053 ( .I(n5760), .ZN(n5739) );
  INVD1BWP U6054 ( .I(n5740), .ZN(n5722) );
  INVD1BWP U6055 ( .I(n5727), .ZN(n5719) );
  INVD1BWP U6056 ( .I(result[6]), .ZN(n4661) );
  ND2D1BWP U6057 ( .A1(\alu/N988 ), .A2(n3925), .ZN(n3851) );
  ND2D1BWP U6058 ( .A1(n5716), .A2(n5715), .ZN(n5720) );
  ND2D1BWP U6059 ( .A1(n4665), .A2(n4668), .ZN(n4059) );
  ND2D1BWP U6060 ( .A1(\alu/N984 ), .A2(n3925), .ZN(n3812) );
  INVD1BWP U6061 ( .I(result[4]), .ZN(n4665) );
  ND2D1BWP U6062 ( .A1(\alu/N986 ), .A2(n3925), .ZN(n3835) );
  INVD1BWP U6063 ( .I(n4672), .ZN(n3913) );
  INVD1BWP U6064 ( .I(n5716), .ZN(n5714) );
  ND2D1BWP U6065 ( .A1(n5708), .A2(n5707), .ZN(n5709) );
  INVD1BWP U6066 ( .I(n4671), .ZN(n3912) );
  INVD1BWP U6067 ( .I(n4690), .ZN(n4054) );
  ND2D1BWP U6068 ( .A1(n4859), .A2(n4701), .ZN(n4861) );
  INVD1BWP U6069 ( .I(n4858), .ZN(n4701) );
  AN2XD1BWP U6070 ( .A1(n4860), .A2(n5616), .Z(n4859) );
  ND2D1BWP U6071 ( .A1(n4862), .A2(op1[1]), .ZN(n4860) );
  ND2D1BWP U6072 ( .A1(n3736), .A2(n3735), .ZN(n3925) );
  INVD1BWP U6073 ( .I(n4691), .ZN(n3735) );
  ND2D1BWP U6074 ( .A1(n3733), .A2(n3734), .ZN(n3739) );
  INVD1BWP U6075 ( .I(n1), .ZN(n3733) );
  INVD1BWP U6076 ( .I(n4692), .ZN(n3736) );
  INVD1BWP U6077 ( .I(func[0]), .ZN(n3734) );
  INVD1BWP U6078 ( .I(n5800), .ZN(n5801) );
  ND2D1BWP U6079 ( .A1(n5795), .A2(n5794), .ZN(n5800) );
  INVD1BWP U6080 ( .I(n5795), .ZN(n5792) );
  ND2D1BWP U6081 ( .A1(n5610), .A2(n5609), .ZN(n5611) );
  INVD1BWP U6082 ( .I(\mult_x_153/n84 ), .ZN(n5799) );
  AN2XD1BWP U6083 ( .A1(n5796), .A2(n5797), .Z(n5798) );
  INVD1BWP U6084 ( .I(\mult_x_153/n79 ), .ZN(n5797) );
  INVD1BWP U6085 ( .I(\mult_x_153/n96 ), .ZN(n5600) );
  INVD1BWP U6086 ( .I(\mult_x_153/n92 ), .ZN(n5601) );
  INVD1BWP U6087 ( .I(\mult_x_153/n102 ), .ZN(n5596) );
  INVD1BWP U6088 ( .I(n5592), .ZN(n5593) );
  INVD1BWP U6089 ( .I(n5588), .ZN(n5594) );
  INVD1BWP U6090 ( .I(n4856), .ZN(n5556) );
  ND2D1BWP U6091 ( .A1(n5606), .A2(n5608), .ZN(n5609) );
  ND2D1BWP U6092 ( .A1(n4689), .A2(n3781), .ZN(n3901) );
  INVD1BWP U6093 ( .I(n5754), .ZN(n3781) );
  ND2D1BWP U6094 ( .A1(n4656), .A2(n5786), .ZN(n5754) );
  INVD1BWP U6095 ( .I(n5756), .ZN(n5761) );
  ND2D1BWP U6096 ( .A1(n4674), .A2(n5705), .ZN(n5724) );
  ND2D1BWP U6097 ( .A1(op2[12]), .A2(n5641), .ZN(n5628) );
  INVD1BWP U6098 ( .I(n3888), .ZN(n3892) );
  INVD1BWP U6099 ( .I(n4645), .ZN(n5706) );
  INVD1BWP U6100 ( .I(n5713), .ZN(n5697) );
  ND2D1BWP U6101 ( .A1(n5698), .A2(n5712), .ZN(n5699) );
  ND2D1BWP U6102 ( .A1(n4441), .A2(n4434), .ZN(n4417) );
  ND2D1BWP U6103 ( .A1(n4453), .A2(n4434), .ZN(n4435) );
  INVD1BWP U6104 ( .I(n4452), .ZN(n4433) );
  INVD1BWP U6105 ( .I(n4414), .ZN(n4437) );
  ND2D1BWP U6106 ( .A1(n4441), .A2(n4454), .ZN(n4442) );
  INVD1BWP U6107 ( .I(n4438), .ZN(n4447) );
  INVD1BWP U6108 ( .I(n4453), .ZN(n4444) );
  ND2D1BWP U6109 ( .A1(n5721), .A2(n4446), .ZN(n4445) );
  ND2D1BWP U6110 ( .A1(n4457), .A2(n4453), .ZN(n3880) );
  INVD1BWP U6111 ( .I(\intadd_35/B[1] ), .ZN(n4419) );
  ND2D1BWP U6112 ( .A1(n4455), .A2(\intadd_35/B[2] ), .ZN(n4448) );
  INVD1BWP U6113 ( .I(\intadd_35/B[0] ), .ZN(n3878) );
  ND2D1BWP U6114 ( .A1(\intadd_35/B[0] ), .A2(n4441), .ZN(n4452) );
  INVD1BWP U6115 ( .I(n5777), .ZN(n5770) );
  INVD1BWP U6116 ( .I(n5779), .ZN(n5780) );
  ND2D1BWP U6117 ( .A1(n4455), .A2(n3867), .ZN(n4411) );
  INVD1BWP U6118 ( .I(n4410), .ZN(n4455) );
  INVD1BWP U6119 ( .I(n4675), .ZN(n3893) );
  INVD1BWP U6120 ( .I(n4456), .ZN(n4423) );
  ND2D1BWP U6121 ( .A1(n4410), .A2(n5693), .ZN(n4413) );
  INVD1BWP U6122 ( .I(n5695), .ZN(n5693) );
  ND2D1BWP U6123 ( .A1(n3870), .A2(n3871), .ZN(n3869) );
  INVD1BWP U6124 ( .I(\intadd_35/A[1] ), .ZN(n3871) );
  ND2D1BWP U6125 ( .A1(\alu/N683 ), .A2(n5632), .ZN(n5704) );
  ND2D1BWP U6126 ( .A1(op1[12]), .A2(n5640), .ZN(n5633) );
  INVD1BWP U6127 ( .I(n4644), .ZN(n5729) );
  INVD1BWP U6128 ( .I(n5711), .ZN(n4674) );
  ND2D1BWP U6129 ( .A1(n3897), .A2(n4460), .ZN(n5711) );
  ND2D1BWP U6130 ( .A1(\alu/N326 ), .A2(n3875), .ZN(n3765) );
  INVD1BWP U6131 ( .I(n3763), .ZN(n3875) );
  INVD1BWP U6132 ( .I(\alu/N337 ), .ZN(n4429) );
  ND2D1BWP U6133 ( .A1(n4458), .A2(n4459), .ZN(n4462) );
  INVD1BWP U6134 ( .I(n3779), .ZN(n4459) );
  ND2D1BWP U6135 ( .A1(n3771), .A2(n3764), .ZN(n3874) );
  INVD1BWP U6136 ( .I(n3798), .ZN(n4425) );
  INVD1BWP U6137 ( .I(\alu/N333 ), .ZN(n3873) );
  INVD1BWP U6138 ( .I(\alu/N330 ), .ZN(n3759) );
  INVD1BWP U6139 ( .I(\alu/N334 ), .ZN(n3872) );
  ND2D1BWP U6140 ( .A1(n3885), .A2(n4428), .ZN(n4410) );
  INVD1BWP U6141 ( .I(\alu/N339 ), .ZN(n3885) );
  INVD1BWP U6142 ( .I(n3894), .ZN(n3884) );
  INVD1BWP U6143 ( .I(\alu/N338 ), .ZN(n4428) );
  ND2D1BWP U6144 ( .A1(n4456), .A2(n3864), .ZN(n3867) );
  INVD1BWP U6145 ( .I(n3772), .ZN(n3866) );
  ND2D1BWP U6146 ( .A1(n3771), .A2(n3770), .ZN(n3865) );
  INVD1BWP U6147 ( .I(\DP_OP_493J11_130_7648/n42 ), .ZN(n3659) );
  INVD1BWP U6148 ( .I(\DP_OP_493J11_130_7648/n13 ), .ZN(n3658) );
  INVD1BWP U6149 ( .I(n3983), .ZN(n4018) );
  INVD1BWP U6150 ( .I(n4752), .ZN(n4019) );
  INVD1BWP U6151 ( .I(n3982), .ZN(n4016) );
  INVD1BWP U6152 ( .I(n4731), .ZN(n4017) );
  INVD1BWP U6153 ( .I(n3987), .ZN(n4024) );
  INVD1BWP U6154 ( .I(n3986), .ZN(n4022) );
  INVD1BWP U6155 ( .I(n3993), .ZN(n4028) );
  INVD1BWP U6156 ( .I(n3992), .ZN(n4027) );
  ND2D1BWP U6157 ( .A1(op2[0]), .A2(n5622), .ZN(n3979) );
  INVD1BWP U6158 ( .I(n4049), .ZN(n4034) );
  ND2D1BWP U6159 ( .A1(op1[0]), .A2(n5622), .ZN(n3978) );
  ND2D1BWP U6160 ( .A1(n5622), .A2(n3652), .ZN(n3988) );
  INVD1BWP U6161 ( .I(n4043), .ZN(n4044) );
  INVD1BWP U6162 ( .I(n3998), .ZN(n4038) );
  INVD1BWP U6163 ( .I(n4735), .ZN(n4051) );
  INVD1BWP U6164 ( .I(n4715), .ZN(n4046) );
  INVD1BWP U6165 ( .I(n4003), .ZN(n4006) );
  INVD1BWP U6166 ( .I(n3969), .ZN(n4040) );
  INVD1BWP U6167 ( .I(n3968), .ZN(n4039) );
  INVD1BWP U6168 ( .I(n4747), .ZN(n4013) );
  INVD1BWP U6169 ( .I(n4727), .ZN(n4011) );
  ND2D1BWP U6170 ( .A1(n4649), .A2(\alu/N87 ), .ZN(n3961) );
  ND2D1BWP U6171 ( .A1(n4649), .A2(\alu/N88 ), .ZN(n3959) );
  INVD1BWP U6172 ( .I(n4008), .ZN(n3955) );
  ND2D1BWP U6173 ( .A1(n3677), .A2(\alu/N88 ), .ZN(n3954) );
  INVD1BWP U6174 ( .I(n4007), .ZN(n3956) );
  ND2D1BWP U6175 ( .A1(n3677), .A2(\alu/N87 ), .ZN(n3953) );
  ND2D1BWP U6176 ( .A1(n3989), .A2(n5692), .ZN(n3957) );
  ND2D1BWP U6177 ( .A1(n4646), .A2(n3678), .ZN(n4715) );
  ND2D1BWP U6178 ( .A1(n4650), .A2(n3989), .ZN(n3958) );
  INVD1BWP U6179 ( .I(n3972), .ZN(n3975) );
  ND2D1BWP U6180 ( .A1(n4647), .A2(n3678), .ZN(n4735) );
  INVD1BWP U6181 ( .I(\alu/N87 ), .ZN(n3964) );
  INVD1BWP U6182 ( .I(\alu/N88 ), .ZN(n3962) );
  ND2D1BWP U6183 ( .A1(n4650), .A2(n3972), .ZN(n3966) );
  ND2D1BWP U6184 ( .A1(n3952), .A2(\alu/N88 ), .ZN(n3969) );
  ND2D1BWP U6185 ( .A1(n3972), .A2(n5692), .ZN(n3967) );
  INVD1BWP U6186 ( .I(\alu/N683 ), .ZN(n4640) );
  INVD1BWP U6187 ( .I(\alu/N684 ), .ZN(n4658) );
  INVD1BWP U6188 ( .I(n4753), .ZN(n3999) );
  INVD1BWP U6189 ( .I(op1[12]), .ZN(n4660) );
  INVD1BWP U6190 ( .I(op2[12]), .ZN(n4077) );
  INVD1BWP U6191 ( .I(n4839), .ZN(n4838) );
  ND2D1BWP U6192 ( .A1(n3952), .A2(\alu/N87 ), .ZN(n3968) );
  ND2D1BWP U6193 ( .A1(n4677), .A2(n4678), .ZN(n5630) );
  INVD1BWP U6194 ( .I(n4751), .ZN(n4649) );
  INVD1BWP U6195 ( .I(op2[11]), .ZN(n4693) );
  ND2D1BWP U6196 ( .A1(op2[11]), .A2(n4678), .ZN(n3949) );
  ND2D1BWP U6197 ( .A1(n3678), .A2(n3677), .ZN(n3960) );
  INVD1BWP U6198 ( .I(n5622), .ZN(n3677) );
  INVD1BWP U6199 ( .I(\intadd_36/B[0] ), .ZN(n3950) );
  INVD1BWP U6200 ( .I(op2[10]), .ZN(n4676) );
  INVD1BWP U6201 ( .I(n3652), .ZN(n3678) );
  INVD1BWP U6202 ( .I(op1[11]), .ZN(n4678) );
  ND2D1BWP U6203 ( .A1(op2[10]), .A2(n4677), .ZN(n5629) );
  INVD1BWP U6204 ( .I(op1[10]), .ZN(n4677) );
  ND2D1BWP U6205 ( .A1(op2[15]), .A2(op1[15]), .ZN(n4056) );
  ND2D1BWP U6206 ( .A1(n3731), .A2(n3730), .ZN(n5240) );
  ND2D1BWP U6207 ( .A1(n3944), .A2(instrIn[11]), .ZN(n3730) );
  INVD1BWP U6208 ( .I(n5200), .ZN(n3731) );
  INVD1BWP U6209 ( .I(n5226), .ZN(n3673) );
  INVD1BWP U6210 ( .I(vectorData2[141]), .ZN(n5216) );
  INVD1BWP U6211 ( .I(n5185), .ZN(n3752) );
  INVD1BWP U6212 ( .I(n5186), .ZN(n3751) );
  INVD1BWP U6213 ( .I(vectorToLoad[195]), .ZN(n6043) );
  INVD1BWP U6214 ( .I(vectorToLoad[194]), .ZN(n6042) );
  INVD1BWP U6215 ( .I(vectorToLoad[193]), .ZN(n6041) );
  ND2D1BWP U6216 ( .A1(n4992), .A2(n4698), .ZN(n4996) );
  ND2D1BWP U6217 ( .A1(cycles[3]), .A2(cycles[2]), .ZN(n4994) );
  ND2D1BWP U6218 ( .A1(n134), .A2(n132), .ZN(n5252) );
  INVD1BWP U6219 ( .I(n3672), .ZN(n3671) );
  INVD1BWP U6220 ( .I(n5213), .ZN(n3672) );
  ND2D1BWP U6221 ( .A1(cycles[2]), .A2(n132), .ZN(n4993) );
  ND2D1BWP U6222 ( .A1(n3745), .A2(n3729), .ZN(n3747) );
  ND2D1BWP U6223 ( .A1(n3728), .A2(n4567), .ZN(n3729) );
  INVD1BWP U6224 ( .I(instrIn[7]), .ZN(n4559) );
  INVD1BWP U6225 ( .I(n3749), .ZN(n3745) );
  INVD1BWP U6226 ( .I(vectorToLoad[223]), .ZN(n6061) );
  INVD1BWP U6227 ( .I(vectorToLoad[222]), .ZN(n6060) );
  INVD1BWP U6228 ( .I(vectorToLoad[220]), .ZN(n6059) );
  INVD1BWP U6229 ( .I(vectorToLoad[219]), .ZN(n6058) );
  INVD1BWP U6230 ( .I(vectorToLoad[218]), .ZN(n6057) );
  INVD1BWP U6231 ( .I(vectorToLoad[217]), .ZN(n6056) );
  INVD1BWP U6232 ( .I(vectorToLoad[216]), .ZN(n6055) );
  INVD1BWP U6233 ( .I(vectorToLoad[215]), .ZN(n6054) );
  INVD1BWP U6234 ( .I(vectorToLoad[214]), .ZN(n6053) );
  INVD1BWP U6235 ( .I(vectorToLoad[212]), .ZN(n6052) );
  INVD1BWP U6236 ( .I(vectorToLoad[211]), .ZN(n6051) );
  INVD1BWP U6237 ( .I(vectorToLoad[209]), .ZN(n6050) );
  INVD1BWP U6238 ( .I(vectorToLoad[207]), .ZN(n6049) );
  INVD1BWP U6239 ( .I(vectorToLoad[205]), .ZN(n6048) );
  INVD1BWP U6240 ( .I(vectorToLoad[204]), .ZN(n6047) );
  INVD1BWP U6241 ( .I(vectorToLoad[203]), .ZN(n6046) );
  INVD1BWP U6242 ( .I(vectorToLoad[201]), .ZN(n6045) );
  INVD1BWP U6243 ( .I(vectorToLoad[197]), .ZN(n6044) );
  ND2D1BWP U6244 ( .A1(op2[0]), .A2(n4815), .ZN(n5587) );
  INVD1BWP U6245 ( .I(n4783), .ZN(\mult_x_153/n94 ) );
  INVD1BWP U6246 ( .I(n4767), .ZN(\mult_x_153/n47 ) );
  INVD1BWP U6247 ( .I(n4844), .ZN(n4845) );
  INVD1BWP U6248 ( .I(n4761), .ZN(\mult_x_153/n42 ) );
  INVD1BWP U6249 ( .I(n4766), .ZN(n4760) );
  INVD1BWP U6250 ( .I(n4769), .ZN(\mult_x_153/n86 ) );
  INVD1BWP U6251 ( .I(n4853), .ZN(n4852) );
  INVD1BWP U6252 ( .I(n4779), .ZN(\mult_x_153/n93 ) );
  INVD1BWP U6253 ( .I(n4849), .ZN(n4801) );
  INVD1BWP U6254 ( .I(n5572), .ZN(n5576) );
  INVD1BWP U6255 ( .I(n6072), .ZN(\mult_x_153/n37 ) );
  INVD1BWP U6256 ( .I(n6071), .ZN(\mult_x_153/n70 ) );
  INVD1BWP U6257 ( .I(op2[2]), .ZN(n4670) );
  INVD1BWP U6258 ( .I(op2[7]), .ZN(n4833) );
  INVD1BWP U6259 ( .I(n5557), .ZN(n5562) );
  ND2D1BWP U6260 ( .A1(op1[3]), .A2(n4669), .ZN(n5566) );
  INVD1BWP U6261 ( .I(op1[2]), .ZN(n4669) );
  ND2D1BWP U6262 ( .A1(op1[2]), .A2(n5561), .ZN(n4768) );
  INVD1BWP U6263 ( .I(op2[3]), .ZN(n5569) );
  INVD1BWP U6264 ( .I(n4817), .ZN(n4816) );
  ND2D1BWP U6265 ( .A1(op1[4]), .A2(n4832), .ZN(n4809) );
  INVD1BWP U6266 ( .I(n4820), .ZN(n4815) );
  ND2D1BWP U6267 ( .A1(n4666), .A2(n5561), .ZN(n5613) );
  INVD1BWP U6268 ( .I(op1[4]), .ZN(n4666) );
  INVD1BWP U6269 ( .I(n4806), .ZN(n4803) );
  ND2D1BWP U6270 ( .A1(op1[6]), .A2(n5605), .ZN(n4798) );
  INVD1BWP U6271 ( .I(n4808), .ZN(n4800) );
  ND2D1BWP U6272 ( .A1(n4662), .A2(n4832), .ZN(n5614) );
  INVD1BWP U6273 ( .I(op1[6]), .ZN(n4662) );
  ND2D1BWP U6274 ( .A1(op2[0]), .A2(n5555), .ZN(n4782) );
  INVD1BWP U6275 ( .I(n4796), .ZN(n4793) );
  INVD1BWP U6276 ( .I(op2[0]), .ZN(n4680) );
  ND2D1BWP U6277 ( .A1(n5612), .A2(n5604), .ZN(n5554) );
  ND2D1BWP U6278 ( .A1(n4653), .A2(n5605), .ZN(n5612) );
  INVD1BWP U6279 ( .I(op1[8]), .ZN(n4653) );
  INVD1BWP U6280 ( .I(op2[6]), .ZN(n4663) );
  INVD1BWP U6281 ( .I(n5573), .ZN(\mult_x_153/n176 ) );
  ND2D1BWP U6282 ( .A1(op1[0]), .A2(op1[1]), .ZN(n5573) );
  INVD1BWP U6283 ( .I(n4827), .ZN(n5570) );
  ND2D1BWP U6284 ( .A1(op1[0]), .A2(n6070), .ZN(n4827) );
  INVD1BWP U6285 ( .I(op1[1]), .ZN(n6070) );
  ND2D1BWP U6286 ( .A1(op1[1]), .A2(n4679), .ZN(n5564) );
  INVD1BWP U6287 ( .I(n4567), .ZN(n4566) );
  NR3D1BWP U6288 ( .A1(\vrf/N12 ), .A2(\vrf/N13 ), .A3(n4622), .ZN(n6080) );
  ND2D1BWP U6289 ( .A1(\vrf/N12 ), .A2(\vrf/N13 ), .ZN(n6078) );
  ND2D1BWP U6290 ( .A1(\vrf/N12 ), .A2(n4620), .ZN(n6076) );
  ND2D1BWP U6291 ( .A1(\vrf/N13 ), .A2(n4621), .ZN(n6074) );
  NR3D1BWP U6292 ( .A1(\vrf/N14 ), .A2(\vrf/N12 ), .A3(\vrf/N13 ), .ZN(n6073)
         );
  INVD1BWP U6293 ( .I(n5985), .ZN(n4562) );
  INVD1BWP U6294 ( .I(n5979), .ZN(n4563) );
  INVD1BWP U6295 ( .I(n5982), .ZN(n4564) );
  ND2D1BWP U6296 ( .A1(n5807), .A2(n137), .ZN(n5814) );
  NR4D1BWP U6297 ( .A1(cycles[4]), .A2(n132), .A3(n5812), .A4(n5811), .ZN(
        n5980) );
  INVD1BWP U6298 ( .I(n134), .ZN(n5817) );
  INVD1BWP U6299 ( .I(n136), .ZN(n5818) );
  ND2D1BWP U6300 ( .A1(cycles[1]), .A2(cycles[2]), .ZN(n5813) );
  ND2D1BWP U6301 ( .A1(cycles[2]), .A2(n136), .ZN(n5810) );
  INVD1BWP U6302 ( .I(n5294), .ZN(n5805) );
  ND2D1BWP U6303 ( .A1(n137), .A2(n5806), .ZN(n5809) );
  ND2D1BWP U6304 ( .A1(n5807), .A2(cycles[0]), .ZN(n5816) );
  ND2D1BWP U6305 ( .A1(cycles[1]), .A2(n134), .ZN(n5808) );
  ND2D1BWP U6306 ( .A1(cycles[0]), .A2(n5806), .ZN(n5815) );
  INVD1BWP U6307 ( .I(\vrf/N14 ), .ZN(n4622) );
  ND2D1BWP U6308 ( .A1(\vrf/N12 ), .A2(\vrf/N13 ), .ZN(n8208) );
  ND2D1BWP U6309 ( .A1(\vrf/N12 ), .A2(n4620), .ZN(n8206) );
  INVD1BWP U6310 ( .I(\vrf/N13 ), .ZN(n4620) );
  ND2D1BWP U6311 ( .A1(\vrf/N13 ), .A2(n4621), .ZN(n8204) );
  INVD1BWP U6312 ( .I(\vrf/N12 ), .ZN(n4621) );
  INVD1BWP U6313 ( .I(instrIn[9]), .ZN(n4557) );
  ND2D1BWP U6314 ( .A1(n3657), .A2(n3656), .ZN(N155) );
  ND2D1BWP U6315 ( .A1(n4542), .A2(n3710), .ZN(n3715) );
  ND2D1BWP U6316 ( .A1(n3727), .A2(n3699), .ZN(n3750) );
  NR3D0BWP U6317 ( .A1(code[2]), .A2(code[3]), .A3(n4697), .ZN(n3727) );
  INVD1BWP U6318 ( .I(n3688), .ZN(n3690) );
  ND2D1BWP U6319 ( .A1(cycles[3]), .A2(n134), .ZN(n4998) );
  ND2D1BWP U6320 ( .A1(n132), .A2(cycles[1]), .ZN(n3685) );
  ND2D1BWP U6321 ( .A1(n3688), .A2(n3728), .ZN(n3686) );
  INVD1BWP U6322 ( .I(n3748), .ZN(n4392) );
  OR3XD1BWP U6323 ( .A1(code[1]), .A2(code[2]), .A3(code[3]), .Z(n3748) );
  ND2D1BWP U6324 ( .A1(n3683), .A2(n4697), .ZN(n3728) );
  INVD1BWP U6325 ( .I(n3786), .ZN(n3683) );
  NR2XD0BWP U6326 ( .A1(n4572), .A2(n4616), .ZN(n4571) );
  ND2D1BWP U6327 ( .A1(n4534), .A2(n4470), .ZN(n3662) );
  NR2XD0BWP U6328 ( .A1(n4994), .A2(n5811), .ZN(n4991) );
  NR2XD0BWP U6329 ( .A1(n4572), .A2(n4068), .ZN(n4574) );
  ND2D1BWP U6330 ( .A1(n4550), .A2(n4399), .ZN(n4401) );
  NR2XD0BWP U6331 ( .A1(n6037), .A2(n5285), .ZN(n5553) );
  NR2XD0BWP U6332 ( .A1(\intadd_34/A[3] ), .A2(n5285), .ZN(n5552) );
  INVD1BWP U6333 ( .I(n4696), .ZN(n3784) );
  NR2XD0BWP U6334 ( .A1(n3679), .A2(n5277), .ZN(n5320) );
  NR2XD0BWP U6335 ( .A1(n3679), .A2(n5278), .ZN(n5322) );
  NR2XD0BWP U6336 ( .A1(n4665), .A2(n5285), .ZN(n5542) );
  NR2XD0BWP U6337 ( .A1(n4664), .A2(n5285), .ZN(n5543) );
  NR2XD0BWP U6338 ( .A1(n4661), .A2(n5285), .ZN(n5544) );
  NR2XD0BWP U6339 ( .A1(n4655), .A2(n5285), .ZN(n5545) );
  NR2XD0BWP U6340 ( .A1(n4652), .A2(n5285), .ZN(n5546) );
  NR2XD0BWP U6341 ( .A1(n4651), .A2(n5285), .ZN(n5547) );
  NR2XD0BWP U6342 ( .A1(n4699), .A2(n5285), .ZN(n5548) );
  NR2XD0BWP U6343 ( .A1(\intadd_34/A[0] ), .A2(n5285), .ZN(n5549) );
  NR2XD0BWP U6344 ( .A1(\intadd_34/A[1] ), .A2(n5285), .ZN(n5550) );
  NR2XD0BWP U6345 ( .A1(n6011), .A2(n5285), .ZN(n5541) );
  NR2XD0BWP U6346 ( .A1(n3679), .A2(n5273), .ZN(n5312) );
  NR2XD0BWP U6347 ( .A1(n4668), .A2(n5285), .ZN(n5540) );
  NR2XD0BWP U6348 ( .A1(n4643), .A2(n5285), .ZN(n5539) );
  NR2XD0BWP U6349 ( .A1(n3679), .A2(n5274), .ZN(n5314) );
  NR2XD0BWP U6350 ( .A1(n3679), .A2(n5275), .ZN(n5316) );
  AN3XD1BWP U6351 ( .A1(n5291), .A2(n5292), .A3(n5290), .Z(n3617) );
  NR2XD0BWP U6352 ( .A1(n3679), .A2(n5281), .ZN(n5328) );
  NR2XD0BWP U6353 ( .A1(n3679), .A2(n5268), .ZN(n5301) );
  NR2XD0BWP U6354 ( .A1(n3679), .A2(n5269), .ZN(n5304) );
  NR2XD0BWP U6355 ( .A1(n3679), .A2(n5276), .ZN(n5318) );
  NR2XD0BWP U6356 ( .A1(n3679), .A2(n5270), .ZN(n5306) );
  AO21D1BWP U6357 ( .A1(n3675), .A2(n5251), .B(n5295), .Z(n4400) );
  NR2XD0BWP U6358 ( .A1(n3679), .A2(n5271), .ZN(n5308) );
  NR2XD0BWP U6359 ( .A1(n3679), .A2(n5272), .ZN(n5310) );
  NR2XD0BWP U6360 ( .A1(\intadd_34/A[2] ), .A2(n5285), .ZN(n5551) );
  ND2D1BWP U6361 ( .A1(cycles[0]), .A2(n5818), .ZN(n5285) );
  INVD1BWP U6362 ( .I(n5368), .ZN(n4547) );
  ND2D1BWP U6363 ( .A1(n5291), .A2(n4990), .ZN(n5368) );
  OAI21D1BWP U6364 ( .A1(n5251), .A2(n3675), .B(n4698), .ZN(n5295) );
  IND2D1BWP U6365 ( .A1(n5298), .B1(n4408), .ZN(n4473) );
  AN2XD1BWP U6366 ( .A1(n5251), .A2(n3675), .Z(n5296) );
  INVD1BWP U6367 ( .I(DataIn[11]), .ZN(n5278) );
  INVD1BWP U6368 ( .I(DataIn[1]), .ZN(n5268) );
  INVD1BWP U6369 ( .I(DataIn[2]), .ZN(n5269) );
  INVD1BWP U6370 ( .I(DataIn[3]), .ZN(n5270) );
  INVD1BWP U6371 ( .I(DataIn[4]), .ZN(n5271) );
  INVD1BWP U6372 ( .I(DataIn[5]), .ZN(n5272) );
  INVD1BWP U6373 ( .I(DataIn[6]), .ZN(n5273) );
  INVD1BWP U6374 ( .I(DataIn[7]), .ZN(n5274) );
  INVD1BWP U6375 ( .I(DataIn[8]), .ZN(n5275) );
  INVD1BWP U6376 ( .I(DataIn[9]), .ZN(n5276) );
  NR2XD0BWP U6377 ( .A1(n4472), .A2(n4471), .ZN(n4477) );
  NR2XD0BWP U6378 ( .A1(n5817), .A2(cycles[1]), .ZN(n5254) );
  NR2XD0BWP U6379 ( .A1(n3788), .A2(n4551), .ZN(n4072) );
  INVD1BWP U6380 ( .I(n4398), .ZN(n4478) );
  INVD1BWP U6381 ( .I(scalarToLoad[15]), .ZN(n4336) );
  INR3D0BWP U6382 ( .A1(n4643), .B1(n4059), .B2(n4058), .ZN(n5247) );
  INVD1BWP U6383 ( .I(result[2]), .ZN(n4668) );
  OAI21D1BWP U6384 ( .A1(func[2]), .A2(func[0]), .B(func[3]), .ZN(n3737) );
  ND2D1BWP U6385 ( .A1(func[2]), .A2(n3733), .ZN(n3738) );
  NR2XD0BWP U6386 ( .A1(n3734), .A2(n3740), .ZN(n4692) );
  NR2XD0BWP U6387 ( .A1(op2[15]), .A2(op1[15]), .ZN(n4055) );
  NR2XD0BWP U6388 ( .A1(n3750), .A2(n3749), .ZN(n4688) );
  NR2XD0BWP U6389 ( .A1(n3747), .A2(n153), .ZN(n5200) );
  NR2XD0BWP U6390 ( .A1(n4542), .A2(n4616), .ZN(n3749) );
  INVD1BWP U6391 ( .I(op2[9]), .ZN(n4648) );
  INVD1BWP U6392 ( .I(op2[8]), .ZN(n4654) );
  INVD1BWP U6393 ( .I(op2[4]), .ZN(n4667) );
  INVD1BWP U6394 ( .I(op2[5]), .ZN(n5615) );
  INVD1BWP U6395 ( .I(op2[1]), .ZN(n5616) );
  INVD1BWP U6396 ( .I(n5554), .ZN(n5555) );
  INVD1BWP U6397 ( .I(op1[0]), .ZN(n4679) );
  ND4D1BWP U6398 ( .A1(WR), .A2(n5828), .A3(n5829), .A4(n4565), .ZN(n4568) );
  INVD1BWP U6399 ( .I(instrIn[10]), .ZN(n4560) );
  INVD1BWP U6400 ( .I(instrIn[11]), .ZN(n4555) );
  ND2D1BWP U6401 ( .A1(n3716), .A2(n3563), .ZN(n3732) );
  NR4D0BWP U6402 ( .A1(code[1]), .A2(code[2]), .A3(code[0]), .A4(n3698), .ZN(
        n3787) );
  OAI21D1BWP U6403 ( .A1(n4573), .A2(n4574), .B(n3020), .ZN(N4170) );
  ND3D1BWP U6404 ( .A1(n4394), .A2(n3681), .A3(n3563), .ZN(n3020) );
  NR2XD0BWP U6405 ( .A1(n4472), .A2(n4478), .ZN(n4396) );
  OAI211D1BWP U6406 ( .A1(n5464), .A2(n3662), .B(n5463), .C(n4535), .ZN(N4426)
         );
  AOI22D1BWP U6407 ( .A1(n3669), .A2(vectorToLoad[208]), .B1(n4625), .B2(n5462), .ZN(n5463) );
  OAI222D1BWP U6408 ( .A1(n6050), .A2(n3670), .B1(n3662), .B2(n5467), .C1(
        n5509), .C2(n5466), .ZN(N4427) );
  NR2XD0BWP U6409 ( .A1(n3675), .A2(n5465), .ZN(n5466) );
  OAI222D1BWP U6410 ( .A1(n6051), .A2(n3670), .B1(n3662), .B2(n5473), .C1(
        n5509), .C2(n5472), .ZN(N4429) );
  NR2XD0BWP U6411 ( .A1(n3675), .A2(n5471), .ZN(n5472) );
  OAI222D1BWP U6412 ( .A1(n6052), .A2(n3670), .B1(n3662), .B2(n5476), .C1(
        n5509), .C2(n5475), .ZN(N4430) );
  NR2XD0BWP U6413 ( .A1(n3675), .A2(n5474), .ZN(n5475) );
  AO222D1BWP U6414 ( .A1(n3624), .A2(n4548), .B1(n5540), .B2(n3667), .C1(n3669), .C2(vectorToLoad[114]), .Z(N4331) );
  OAI211D1BWP U6415 ( .A1(n5479), .A2(n3662), .B(n5478), .C(n4535), .ZN(N4431)
         );
  AOI22D1BWP U6416 ( .A1(n3669), .A2(vectorToLoad[213]), .B1(n4627), .B2(n5477), .ZN(n5478) );
  OAI211D1BWP U6417 ( .A1(n5470), .A2(n3662), .B(n5469), .C(n4535), .ZN(N4428)
         );
  AOI22D1BWP U6418 ( .A1(n3669), .A2(vectorToLoad[210]), .B1(n4627), .B2(n5468), .ZN(n5469) );
  OAI22D1BWP U6419 ( .A1(n4652), .A2(n5249), .B1(n4906), .B2(n4932), .ZN(N1818) );
  OAI222D1BWP U6420 ( .A1(n6053), .A2(n3670), .B1(n3662), .B2(n5482), .C1(
        n5509), .C2(n5481), .ZN(N4433) );
  NR2XD0BWP U6421 ( .A1(n3675), .A2(n5480), .ZN(n5481) );
  OAI21D1BWP U6422 ( .A1(n4401), .A2(\intadd_34/A[2] ), .B(n5264), .ZN(N4246)
         );
  AOI22D1BWP U6423 ( .A1(n3669), .A2(vectorToLoad[29]), .B1(n4629), .B2(n5408), 
        .ZN(n5264) );
  OAI21D1BWP U6424 ( .A1(\intadd_34/A[3] ), .A2(n4401), .B(n5265), .ZN(N4247)
         );
  AOI22D1BWP U6425 ( .A1(n3669), .A2(vectorToLoad[30]), .B1(n4629), .B2(n5410), 
        .ZN(n5265) );
  AO222D1BWP U6426 ( .A1(n3623), .A2(n4548), .B1(n5549), .B2(n4628), .C1(n3668), .C2(vectorToLoad[123]), .Z(N4341) );
  OAI222D1BWP U6427 ( .A1(n6054), .A2(n3670), .B1(n3662), .B2(n5485), .C1(
        n5509), .C2(n5484), .ZN(N4434) );
  NR2XD0BWP U6428 ( .A1(n3675), .A2(n5483), .ZN(n5484) );
  OAI21D1BWP U6429 ( .A1(n4401), .A2(n6037), .B(n5266), .ZN(N4248) );
  AOI22D1BWP U6430 ( .A1(n3669), .A2(vectorToLoad[31]), .B1(n4629), .B2(n5412), 
        .ZN(n5266) );
  OAI22D1BWP U6431 ( .A1(n4655), .A2(n5249), .B1(n4931), .B2(n4906), .ZN(N1817) );
  OAI222D1BWP U6432 ( .A1(n6055), .A2(n3670), .B1(n3662), .B2(n5488), .C1(
        n5509), .C2(n5487), .ZN(N4435) );
  NR2XD0BWP U6433 ( .A1(n3675), .A2(n5486), .ZN(n5487) );
  OAI222D1BWP U6434 ( .A1(n6056), .A2(n3670), .B1(n3662), .B2(n5491), .C1(
        n5509), .C2(n5490), .ZN(N4436) );
  NR2XD0BWP U6435 ( .A1(n3675), .A2(n5489), .ZN(n5490) );
  OAI21D1BWP U6436 ( .A1(n4401), .A2(\intadd_34/A[1] ), .B(n5263), .ZN(N4245)
         );
  AOI22D1BWP U6437 ( .A1(n3669), .A2(vectorToLoad[28]), .B1(n4629), .B2(n5406), 
        .ZN(n5263) );
  OAI222D1BWP U6438 ( .A1(n6057), .A2(n3670), .B1(n3662), .B2(n5494), .C1(
        n5509), .C2(n5493), .ZN(N4437) );
  NR2XD0BWP U6439 ( .A1(n3675), .A2(n5492), .ZN(n5493) );
  OAI222D1BWP U6440 ( .A1(n6058), .A2(n3670), .B1(n3662), .B2(n5497), .C1(
        n5509), .C2(n5496), .ZN(N4438) );
  NR2XD0BWP U6441 ( .A1(n3675), .A2(n5495), .ZN(n5496) );
  AO222D1BWP U6442 ( .A1(n3625), .A2(n4548), .B1(n5541), .B2(n3667), .C1(n3668), .C2(vectorToLoad[115]), .Z(N4333) );
  AO222D1BWP U6443 ( .A1(n3633), .A2(n4548), .B1(n5552), .B2(n3667), .C1(n3669), .C2(vectorToLoad[126]), .Z(N4344) );
  OAI222D1BWP U6444 ( .A1(n6059), .A2(n3670), .B1(n3662), .B2(n5500), .C1(
        n5509), .C2(n5499), .ZN(N4439) );
  NR2XD0BWP U6445 ( .A1(n3675), .A2(n5498), .ZN(n5499) );
  AO222D1BWP U6446 ( .A1(n4550), .A2(n5358), .B1(n5357), .B2(n4629), .C1(
        vectorToLoad[27]), .C2(n3668), .Z(N4244) );
  OAI211D1BWP U6447 ( .A1(n5503), .A2(n3662), .B(n5502), .C(n4535), .ZN(N4440)
         );
  AOI22D1BWP U6448 ( .A1(n3669), .A2(vectorToLoad[221]), .B1(n4627), .B2(n5501), .ZN(n5502) );
  OAI22D1BWP U6449 ( .A1(n4906), .A2(n4928), .B1(n4661), .B2(n5249), .ZN(N1816) );
  OAI222D1BWP U6450 ( .A1(n6060), .A2(n3670), .B1(n3662), .B2(n5506), .C1(
        n5509), .C2(n5505), .ZN(N4441) );
  NR2XD0BWP U6451 ( .A1(n3675), .A2(n5504), .ZN(n5505) );
  OAI222D1BWP U6452 ( .A1(n6061), .A2(n3670), .B1(n3662), .B2(n5510), .C1(
        n5509), .C2(n5508), .ZN(N4442) );
  NR2XD0BWP U6453 ( .A1(n3675), .A2(n5507), .ZN(n5508) );
  OAI21D1BWP U6454 ( .A1(n4401), .A2(n4699), .B(n5262), .ZN(N4243) );
  AOI22D1BWP U6455 ( .A1(n3669), .A2(vectorToLoad[26]), .B1(n4629), .B2(n5403), 
        .ZN(n5262) );
  AO211D1BWP U6456 ( .A1(n3668), .A2(vectorToLoad[224]), .B(n4505), .C(n4479), 
        .Z(N4443) );
  AO222D1BWP U6457 ( .A1(n3620), .A2(n4548), .B1(n5539), .B2(n3667), .C1(n3669), .C2(vectorToLoad[113]), .Z(N4330) );
  OAI211D1BWP U6458 ( .A1(n5506), .A2(n4407), .B(n5411), .C(n4535), .ZN(N4408)
         );
  AOI22D1BWP U6459 ( .A1(n3669), .A2(vectorToLoad[190]), .B1(n5415), .B2(n5552), .ZN(n5411) );
  AO222D1BWP U6460 ( .A1(n3648), .A2(n4548), .B1(n5534), .B2(n4628), .C1(n4631), .C2(vectorToLoad[110]), .Z(N4327) );
  OAI211D1BWP U6461 ( .A1(n5510), .A2(n4407), .B(n5413), .C(n4535), .ZN(N4409)
         );
  AOI22D1BWP U6462 ( .A1(n3669), .A2(vectorToLoad[191]), .B1(n5415), .B2(n5553), .ZN(n5413) );
  AO222D1BWP U6463 ( .A1(n3669), .A2(vectorToLoad[36]), .B1(n4549), .B2(n5524), 
        .C1(n3649), .C2(n5308), .Z(N4253) );
  OAI222D1BWP U6464 ( .A1(n6041), .A2(n3670), .B1(n3662), .B2(n5517), .C1(
        n5509), .C2(n5421), .ZN(N4411) );
  NR2XD0BWP U6465 ( .A1(n3675), .A2(n5420), .ZN(n5421) );
  AO222D1BWP U6466 ( .A1(n3631), .A2(n4548), .B1(n5550), .B2(n3667), .C1(n3668), .C2(vectorToLoad[124]), .Z(N4342) );
  OAI222D1BWP U6467 ( .A1(n6042), .A2(n3670), .B1(n3662), .B2(n5520), .C1(
        n5509), .C2(n5423), .ZN(N4412) );
  NR2XD0BWP U6468 ( .A1(n3675), .A2(n5422), .ZN(n5423) );
  OAI222D1BWP U6469 ( .A1(n6043), .A2(n3670), .B1(n3662), .B2(n5523), .C1(
        n5509), .C2(n5425), .ZN(N4413) );
  NR2XD0BWP U6470 ( .A1(n3675), .A2(n5424), .ZN(n5425) );
  AO222D1BWP U6471 ( .A1(n3669), .A2(vectorToLoad[35]), .B1(n5306), .B2(n3649), 
        .C1(n4549), .C2(n5521), .Z(N4252) );
  OAI211D1BWP U6472 ( .A1(n5428), .A2(n3662), .B(n5427), .C(n4535), .ZN(N4414)
         );
  AOI22D1BWP U6473 ( .A1(n3669), .A2(vectorToLoad[196]), .B1(n4627), .B2(n5426), .ZN(n5427) );
  AO222D1BWP U6474 ( .A1(n3636), .A2(n4548), .B1(n5535), .B2(n3667), .C1(n3669), .C2(vectorToLoad[111]), .Z(N4328) );
  OAI222D1BWP U6475 ( .A1(n6044), .A2(n3670), .B1(n3662), .B2(n5431), .C1(
        n5509), .C2(n5430), .ZN(N4415) );
  NR2XD0BWP U6476 ( .A1(n3675), .A2(n5429), .ZN(n5430) );
  OAI211D1BWP U6477 ( .A1(n5434), .A2(n3662), .B(n5433), .C(n4535), .ZN(N4416)
         );
  AOI22D1BWP U6478 ( .A1(n3669), .A2(vectorToLoad[198]), .B1(n4627), .B2(n5432), .ZN(n5433) );
  AO222D1BWP U6479 ( .A1(n3668), .A2(vectorToLoad[34]), .B1(n5304), .B2(n3649), 
        .C1(n4549), .C2(n5518), .Z(N4251) );
  OAI211D1BWP U6480 ( .A1(n5437), .A2(n3662), .B(n5436), .C(n4535), .ZN(N4417)
         );
  AOI22D1BWP U6481 ( .A1(n3669), .A2(vectorToLoad[199]), .B1(n4627), .B2(n5435), .ZN(n5436) );
  OAI211D1BWP U6482 ( .A1(n5440), .A2(n3662), .B(n5439), .C(n4535), .ZN(N4418)
         );
  AOI22D1BWP U6483 ( .A1(n3669), .A2(vectorToLoad[200]), .B1(n4627), .B2(n5438), .ZN(n5439) );
  OAI222D1BWP U6484 ( .A1(n6045), .A2(n3670), .B1(n3662), .B2(n5443), .C1(
        n5509), .C2(n5442), .ZN(N4419) );
  NR2XD0BWP U6485 ( .A1(n3675), .A2(n5441), .ZN(n5442) );
  AO222D1BWP U6486 ( .A1(n3668), .A2(vectorToLoad[33]), .B1(n5301), .B2(n3649), 
        .C1(n4549), .C2(n5515), .Z(N4250) );
  OAI211D1BWP U6487 ( .A1(n5446), .A2(n3662), .B(n5445), .C(n4535), .ZN(N4420)
         );
  AOI22D1BWP U6488 ( .A1(n3669), .A2(vectorToLoad[202]), .B1(n4627), .B2(n5444), .ZN(n5445) );
  AO222D1BWP U6489 ( .A1(n3668), .A2(vectorToLoad[112]), .B1(n3667), .B2(n5536), .C1(n4548), .C2(n5537), .Z(N4329) );
  OAI222D1BWP U6490 ( .A1(n6046), .A2(n3670), .B1(n3662), .B2(n5449), .C1(
        n5509), .C2(n5448), .ZN(N4421) );
  NR2XD0BWP U6491 ( .A1(n3675), .A2(n5447), .ZN(n5448) );
  OAI222D1BWP U6492 ( .A1(n6047), .A2(n3670), .B1(n3662), .B2(n5452), .C1(
        n5509), .C2(n5451), .ZN(N4422) );
  NR2XD0BWP U6493 ( .A1(n3675), .A2(n5450), .ZN(n5451) );
  OAI22D1BWP U6494 ( .A1(n4651), .A2(n5249), .B1(n4961), .B2(n4909), .ZN(N1819) );
  AO222D1BWP U6495 ( .A1(n3668), .A2(vectorToLoad[32]), .B1(n4549), .B2(n5511), 
        .C1(n3649), .C2(n5297), .Z(N4249) );
  OAI222D1BWP U6496 ( .A1(n6048), .A2(n3670), .B1(n3662), .B2(n5455), .C1(
        n5509), .C2(n5454), .ZN(N4423) );
  NR2XD0BWP U6497 ( .A1(n3675), .A2(n5453), .ZN(n5454) );
  AO222D1BWP U6498 ( .A1(n3632), .A2(n4548), .B1(n5551), .B2(n3667), .C1(n4631), .C2(vectorToLoad[125]), .Z(N4343) );
  OAI211D1BWP U6499 ( .A1(n5458), .A2(n3662), .B(n5457), .C(n4535), .ZN(N4424)
         );
  AOI22D1BWP U6500 ( .A1(n3669), .A2(vectorToLoad[206]), .B1(n4627), .B2(n5456), .ZN(n5457) );
  OAI222D1BWP U6501 ( .A1(n6049), .A2(n3670), .B1(n3662), .B2(n5461), .C1(
        n5509), .C2(n5460), .ZN(N4425) );
  NR2XD0BWP U6502 ( .A1(n3675), .A2(n5459), .ZN(n5460) );
  OAI211D1BWP U6503 ( .A1(n3670), .A2(n4515), .B(n4514), .C(n4535), .ZN(N4464)
         );
  AOI22D1BWP U6504 ( .A1(n3665), .A2(n5543), .B1(n4534), .B2(n3626), .ZN(n4514) );
  OAI211D1BWP U6505 ( .A1(n3670), .A2(n4517), .B(n4516), .C(n4535), .ZN(N4465)
         );
  AOI22D1BWP U6506 ( .A1(n3665), .A2(n5544), .B1(n4534), .B2(n3627), .ZN(n4516) );
  OAI211D1BWP U6507 ( .A1(n3670), .A2(n4519), .B(n4518), .C(n4535), .ZN(N4466)
         );
  AOI22D1BWP U6508 ( .A1(n3665), .A2(n5545), .B1(n4534), .B2(n3628), .ZN(n4518) );
  AO222D1BWP U6509 ( .A1(n4550), .A2(n5342), .B1(n5341), .B2(n4629), .C1(
        vectorToLoad[20]), .C2(n3669), .Z(N4237) );
  OAI211D1BWP U6510 ( .A1(n3670), .A2(n4521), .B(n4520), .C(n4535), .ZN(N4467)
         );
  AOI22D1BWP U6511 ( .A1(n3665), .A2(n5546), .B1(n4534), .B2(n3629), .ZN(n4520) );
  OAI211D1BWP U6512 ( .A1(n3670), .A2(n4523), .B(n4522), .C(n4535), .ZN(N4468)
         );
  AOI22D1BWP U6513 ( .A1(n3665), .A2(n5547), .B1(n4534), .B2(n3622), .ZN(n4522) );
  AO222D1BWP U6514 ( .A1(n3630), .A2(n4548), .B1(n5548), .B2(n4628), .C1(n3669), .C2(vectorToLoad[122]), .Z(N4340) );
  OAI211D1BWP U6515 ( .A1(n3670), .A2(n4525), .B(n4524), .C(n4535), .ZN(N4469)
         );
  AOI22D1BWP U6516 ( .A1(n3665), .A2(n5548), .B1(n4534), .B2(n3630), .ZN(n4524) );
  OAI211D1BWP U6517 ( .A1(n3670), .A2(n4527), .B(n4526), .C(n4535), .ZN(N4470)
         );
  AOI22D1BWP U6518 ( .A1(n3665), .A2(n5549), .B1(n4534), .B2(n3623), .ZN(n4526) );
  OAI211D1BWP U6519 ( .A1(n3670), .A2(n4529), .B(n4528), .C(n4535), .ZN(N4471)
         );
  AOI22D1BWP U6520 ( .A1(n3665), .A2(n5550), .B1(n4534), .B2(n3631), .ZN(n4528) );
  OAI211D1BWP U6521 ( .A1(n3670), .A2(n4531), .B(n4530), .C(n4535), .ZN(N4472)
         );
  AOI22D1BWP U6522 ( .A1(n3665), .A2(n5551), .B1(n4534), .B2(n3632), .ZN(n4530) );
  OAI211D1BWP U6523 ( .A1(n3670), .A2(n4533), .B(n4532), .C(n4535), .ZN(N4473)
         );
  AOI22D1BWP U6524 ( .A1(n3665), .A2(n5552), .B1(n4534), .B2(n3633), .ZN(n4532) );
  OAI211D1BWP U6525 ( .A1(n3670), .A2(n4537), .B(n4536), .C(n4535), .ZN(N4474)
         );
  AOI22D1BWP U6526 ( .A1(n3665), .A2(n5553), .B1(n4534), .B2(n3634), .ZN(n4536) );
  OAI21D1BWP U6527 ( .A1(n6011), .A2(n4401), .B(n5257), .ZN(N4236) );
  AOI22D1BWP U6528 ( .A1(n3669), .A2(vectorToLoad[19]), .B1(n4629), .B2(n5391), 
        .ZN(n5257) );
  AO222D1BWP U6529 ( .A1(n3629), .A2(n4548), .B1(n5546), .B2(n3667), .C1(n3668), .C2(vectorToLoad[120]), .Z(N4338) );
  AOI21D1BWP U6530 ( .A1(n5368), .A2(n5419), .B(n4574), .ZN(N4173) );
  OAI22D1BWP U6531 ( .A1(n5249), .A2(n4643), .B1(n4906), .B2(n4913), .ZN(N1811) );
  NR2XD0BWP U6532 ( .A1(n4574), .A2(n4990), .ZN(N4172) );
  NR2XD0BWP U6533 ( .A1(n4574), .A2(cycles[0]), .ZN(N4171) );
  OAI22D1BWP U6534 ( .A1(nextInstrAddr[0]), .A2(n4064), .B1(n6004), .B2(n3939), 
        .ZN(N4153) );
  OAI211D1BWP U6535 ( .A1(n3670), .A2(n4513), .B(n4512), .C(n4535), .ZN(N4463)
         );
  AOI22D1BWP U6536 ( .A1(n3665), .A2(n5542), .B1(n4534), .B2(n3621), .ZN(n4512) );
  OAI31D1BWP U6537 ( .A1(n3838), .A2(n3816), .A3(n4064), .B(n3815), .ZN(N4155)
         );
  AOI21D1BWP U6538 ( .A1(nextInstrAddr[1]), .A2(nextInstrAddr[0]), .B(
        nextInstrAddr[2]), .ZN(n3816) );
  OAI22D1BWP U6539 ( .A1(n6011), .A2(n3939), .B1(n4064), .B2(n3826), .ZN(N4156) );
  XNR2D1BWP U6540 ( .A1(n3838), .A2(nextInstrAddr[3]), .ZN(n3826) );
  OAI21D1BWP U6541 ( .A1(n4668), .A2(n4401), .B(n5256), .ZN(N4235) );
  AOI22D1BWP U6542 ( .A1(n3669), .A2(vectorToLoad[18]), .B1(n4629), .B2(n5389), 
        .ZN(n5256) );
  AO21D1BWP U6543 ( .A1(n4066), .A2(result[4]), .B(n3840), .Z(N4157) );
  OAI31D1BWP U6544 ( .A1(n3858), .A2(n3839), .A3(n4064), .B(n5998), .ZN(n3840)
         );
  AOI21D1BWP U6545 ( .A1(nextInstrAddr[3]), .A2(n3838), .B(nextInstrAddr[4]), 
        .ZN(n3839) );
  OAI211D1BWP U6546 ( .A1(n4064), .A2(n3849), .B(n5998), .C(n3848), .ZN(N4158)
         );
  XNR2D1BWP U6547 ( .A1(n3858), .A2(nextInstrAddr[5]), .ZN(n3849) );
  AO21D1BWP U6548 ( .A1(n4066), .A2(result[6]), .B(n3860), .Z(N4159) );
  OAI31D1BWP U6549 ( .A1(n3922), .A2(n3859), .A3(n4064), .B(n5998), .ZN(n3860)
         );
  AOI21D1BWP U6550 ( .A1(nextInstrAddr[5]), .A2(n3858), .B(nextInstrAddr[6]), 
        .ZN(n3859) );
  OAI211D1BWP U6551 ( .A1(n4064), .A2(n3908), .B(n5998), .C(n3907), .ZN(N4160)
         );
  XNR2D1BWP U6552 ( .A1(nextInstrAddr[7]), .A2(n3922), .ZN(n3908) );
  AO21D1BWP U6553 ( .A1(n4066), .A2(result[8]), .B(n3924), .Z(N4161) );
  OAI31D1BWP U6554 ( .A1(n3929), .A2(n3923), .A3(n4064), .B(n5998), .ZN(n3924)
         );
  AOI21D1BWP U6555 ( .A1(nextInstrAddr[7]), .A2(n3922), .B(nextInstrAddr[8]), 
        .ZN(n3923) );
  OAI22D1BWP U6556 ( .A1(n5249), .A2(n6004), .B1(n4906), .B2(n4937), .ZN(N1810) );
  NR2XD0BWP U6557 ( .A1(n4063), .A2(n4062), .ZN(n4641) );
  OAI211D1BWP U6558 ( .A1(n4064), .A2(n3936), .B(n5998), .C(n3935), .ZN(N4167)
         );
  XOR2D1BWP U6559 ( .A1(nextInstrAddr[13]), .A2(n4062), .Z(n3936) );
  OAI211D1BWP U6560 ( .A1(n4546), .A2(n3670), .B(n4545), .C(n4544), .ZN(N4233)
         );
  NR2XD0BWP U6561 ( .A1(n4540), .A2(n5464), .ZN(n4541) );
  ND3D1BWP U6562 ( .A1(n3932), .A2(nextInstrAddr[11]), .A3(nextInstrAddr[12]), 
        .ZN(n4062) );
  OAI211D1BWP U6563 ( .A1(n4064), .A2(n3934), .B(n5998), .C(n3933), .ZN(N4165)
         );
  XNR2D1BWP U6564 ( .A1(n3932), .A2(nextInstrAddr[11]), .ZN(n3934) );
  OAI21D1BWP U6565 ( .A1(n4643), .A2(n4401), .B(n5255), .ZN(N4234) );
  AOI22D1BWP U6566 ( .A1(n3669), .A2(vectorToLoad[17]), .B1(n4629), .B2(n5387), 
        .ZN(n5255) );
  OAI31D1BWP U6567 ( .A1(n3932), .A2(n3795), .A3(n4064), .B(n3794), .ZN(N4164)
         );
  AOI21D1BWP U6568 ( .A1(n4066), .A2(result[10]), .B(n4065), .ZN(n3794) );
  AOI21D1BWP U6569 ( .A1(n3929), .A2(nextInstrAddr[9]), .B(nextInstrAddr[10]), 
        .ZN(n3795) );
  AO222D1BWP U6570 ( .A1(n3622), .A2(n4548), .B1(n5547), .B2(n3667), .C1(n4631), .C2(vectorToLoad[121]), .Z(N4339) );
  OAI211D1BWP U6571 ( .A1(n4064), .A2(n3931), .B(n5998), .C(n3930), .ZN(N4163)
         );
  XNR2D1BWP U6572 ( .A1(nextInstrAddr[9]), .A2(n3929), .ZN(n3931) );
  NR2XD0BWP U6573 ( .A1(n3806), .A2(Reset), .ZN(n3805) );
  AO222D1BWP U6574 ( .A1(n3621), .A2(n4548), .B1(n5542), .B2(n3667), .C1(n3669), .C2(vectorToLoad[116]), .Z(N4334) );
  OAI211D1BWP U6575 ( .A1(n5517), .A2(n4409), .B(n5516), .C(n4535), .ZN(N4444)
         );
  AOI22D1BWP U6576 ( .A1(n3669), .A2(vectorToLoad[225]), .B1(n4625), .B2(n5515), .ZN(n5516) );
  OAI22D1BWP U6577 ( .A1(n4906), .A2(n4914), .B1(n4664), .B2(n5249), .ZN(N1815) );
  OAI211D1BWP U6578 ( .A1(n5520), .A2(n4409), .B(n5519), .C(n4535), .ZN(N4445)
         );
  AOI22D1BWP U6579 ( .A1(n3669), .A2(vectorToLoad[226]), .B1(n4625), .B2(n5518), .ZN(n5519) );
  AO222D1BWP U6580 ( .A1(n4550), .A2(n5353), .B1(n5352), .B2(n4629), .C1(
        vectorToLoad[25]), .C2(n3668), .Z(N4242) );
  OAI211D1BWP U6581 ( .A1(n5523), .A2(n4409), .B(n5522), .C(n4535), .ZN(N4446)
         );
  AOI22D1BWP U6582 ( .A1(n3669), .A2(vectorToLoad[227]), .B1(n4625), .B2(n5521), .ZN(n5522) );
  OAI211D1BWP U6583 ( .A1(n3670), .A2(n4481), .B(n4480), .C(n4535), .ZN(N4447)
         );
  AOI22D1BWP U6584 ( .A1(n4625), .A2(n5524), .B1(n4534), .B2(n3635), .ZN(n4480) );
  AO222D1BWP U6585 ( .A1(n3626), .A2(n4548), .B1(n5543), .B2(n3667), .C1(n3668), .C2(vectorToLoad[117]), .Z(N4335) );
  OAI211D1BWP U6586 ( .A1(n3670), .A2(n4483), .B(n4482), .C(n4535), .ZN(N4448)
         );
  AOI22D1BWP U6587 ( .A1(n4625), .A2(n5525), .B1(n4534), .B2(n3639), .ZN(n4482) );
  OAI21D1BWP U6588 ( .A1(n4652), .A2(n4401), .B(n5261), .ZN(N4241) );
  AOI22D1BWP U6589 ( .A1(n3669), .A2(vectorToLoad[24]), .B1(n4629), .B2(n5400), 
        .ZN(n5261) );
  OAI211D1BWP U6590 ( .A1(n3670), .A2(n4485), .B(n4484), .C(n4535), .ZN(N4449)
         );
  AOI22D1BWP U6591 ( .A1(n3665), .A2(n5526), .B1(n4534), .B2(n3640), .ZN(n4484) );
  OAI211D1BWP U6592 ( .A1(n3670), .A2(n4487), .B(n4486), .C(n4535), .ZN(N4450)
         );
  AOI22D1BWP U6593 ( .A1(n3665), .A2(n5527), .B1(n4534), .B2(n3641), .ZN(n4486) );
  OAI211D1BWP U6594 ( .A1(n3670), .A2(n4489), .B(n4488), .C(n4535), .ZN(N4451)
         );
  AOI22D1BWP U6595 ( .A1(n3665), .A2(n5528), .B1(n4534), .B2(n3642), .ZN(n4488) );
  OAI22D1BWP U6596 ( .A1(n4906), .A2(n4911), .B1(n5249), .B2(n4665), .ZN(N1814) );
  OAI211D1BWP U6597 ( .A1(n3670), .A2(n4491), .B(n4490), .C(n4535), .ZN(N4452)
         );
  AOI22D1BWP U6598 ( .A1(n3665), .A2(n5529), .B1(n4534), .B2(n3643), .ZN(n4490) );
  OAI21D1BWP U6599 ( .A1(n4655), .A2(n4401), .B(n5260), .ZN(N4240) );
  AOI22D1BWP U6600 ( .A1(n3669), .A2(vectorToLoad[23]), .B1(n4629), .B2(n5398), 
        .ZN(n5260) );
  OAI211D1BWP U6601 ( .A1(n3670), .A2(n4493), .B(n4492), .C(n4535), .ZN(N4453)
         );
  AOI22D1BWP U6602 ( .A1(n3665), .A2(n5530), .B1(n4534), .B2(n3644), .ZN(n4492) );
  OAI211D1BWP U6603 ( .A1(n3670), .A2(n4495), .B(n4494), .C(n4535), .ZN(N4454)
         );
  AOI22D1BWP U6604 ( .A1(n3665), .A2(n5531), .B1(n4534), .B2(n3645), .ZN(n4494) );
  AO222D1BWP U6605 ( .A1(n3627), .A2(n4548), .B1(n5544), .B2(n3667), .C1(n3668), .C2(vectorToLoad[118]), .Z(N4336) );
  OAI211D1BWP U6606 ( .A1(n3670), .A2(n4497), .B(n4496), .C(n4535), .ZN(N4455)
         );
  AOI22D1BWP U6607 ( .A1(n3665), .A2(n5532), .B1(n4534), .B2(n3646), .ZN(n4496) );
  OAI21D1BWP U6608 ( .A1(n4661), .A2(n4401), .B(n5259), .ZN(N4239) );
  AOI22D1BWP U6609 ( .A1(n3669), .A2(vectorToLoad[22]), .B1(n4629), .B2(n5396), 
        .ZN(n5259) );
  OAI22D1BWP U6610 ( .A1(n4906), .A2(n4930), .B1(n5249), .B2(n6011), .ZN(N1813) );
  OAI211D1BWP U6611 ( .A1(n3670), .A2(n4499), .B(n4498), .C(n4535), .ZN(N4456)
         );
  AOI22D1BWP U6612 ( .A1(n3665), .A2(n5533), .B1(n4534), .B2(n3647), .ZN(n4498) );
  OAI211D1BWP U6613 ( .A1(n3670), .A2(n4501), .B(n4500), .C(n4535), .ZN(N4457)
         );
  AOI22D1BWP U6614 ( .A1(n3665), .A2(n5534), .B1(n4534), .B2(n3648), .ZN(n4500) );
  OAI211D1BWP U6615 ( .A1(n3670), .A2(n4503), .B(n4502), .C(n4535), .ZN(N4458)
         );
  AOI22D1BWP U6616 ( .A1(n3665), .A2(n5535), .B1(n4534), .B2(n3636), .ZN(n4502) );
  OAI21D1BWP U6617 ( .A1(n4664), .A2(n4401), .B(n5258), .ZN(N4238) );
  AOI22D1BWP U6618 ( .A1(n3669), .A2(vectorToLoad[21]), .B1(n4629), .B2(n5394), 
        .ZN(n5258) );
  AO211D1BWP U6619 ( .A1(n3668), .A2(vectorToLoad[240]), .B(n4505), .C(n4504), 
        .Z(N4459) );
  NR2XD0BWP U6620 ( .A1(n5805), .A2(n5464), .ZN(n5537) );
  AO222D1BWP U6621 ( .A1(n3634), .A2(n4548), .B1(n5553), .B2(n3667), .C1(n4631), .C2(vectorToLoad[127]), .Z(N4345) );
  OAI211D1BWP U6622 ( .A1(n3670), .A2(n4507), .B(n4506), .C(n4535), .ZN(N4460)
         );
  AOI22D1BWP U6623 ( .A1(n3665), .A2(n5539), .B1(n4534), .B2(n3620), .ZN(n4506) );
  AO222D1BWP U6624 ( .A1(n3628), .A2(n4548), .B1(n5545), .B2(n3667), .C1(n4631), .C2(vectorToLoad[119]), .Z(N4337) );
  OAI211D1BWP U6625 ( .A1(n3670), .A2(n4509), .B(n4508), .C(n4535), .ZN(N4461)
         );
  AOI22D1BWP U6626 ( .A1(n3665), .A2(n5540), .B1(n4534), .B2(n3624), .ZN(n4508) );
  OAI22D1BWP U6627 ( .A1(n5249), .A2(n4668), .B1(n4906), .B2(n4910), .ZN(N1812) );
  OAI211D1BWP U6628 ( .A1(n3670), .A2(n4511), .B(n4510), .C(n4535), .ZN(N4462)
         );
  AOI22D1BWP U6629 ( .A1(n3665), .A2(n5541), .B1(n4534), .B2(n3625), .ZN(n4510) );
  MUX2ND0BWP U6630 ( .I0(n6037), .I1(n4336), .S(n4084), .ZN(N1825) );
  NR2XD0BWP U6631 ( .A1(n3676), .A2(n4474), .ZN(n4084) );
  OAI21D1BWP U6632 ( .A1(n4467), .A2(n4555), .B(n4466), .ZN(N4214) );
  AO222D1BWP U6633 ( .A1(n4550), .A2(n5498), .B1(n3650), .B2(n5406), .C1(
        vectorToLoad[92]), .C2(n4631), .Z(N4309) );
  NR2XD0BWP U6634 ( .A1(n5290), .A2(\intadd_34/A[1] ), .ZN(n5498) );
  AO222D1BWP U6635 ( .A1(n3669), .A2(vectorToLoad[59]), .B1(n5357), .B2(n3649), 
        .C1(n4549), .C2(n5549), .Z(N4276) );
  OAI211D1BWP U6636 ( .A1(n3797), .A2(n4560), .B(n5199), .C(n3796), .ZN(N4202)
         );
  AOI211XD0BWP U6637 ( .A1(n4681), .A2(vectorData2[10]), .B(n5200), .C(n5198), 
        .ZN(n5199) );
  AOI31D1BWP U6638 ( .A1(n5196), .A2(n5195), .A3(n5197), .B(n3661), .ZN(n5198)
         );
  AOI22D1BWP U6639 ( .A1(vectorData2[26]), .A2(n5184), .B1(vectorData2[122]), 
        .B2(n5231), .ZN(n5197) );
  AOI211XD0BWP U6640 ( .A1(vectorData2[218]), .A2(n5228), .B(n5194), .C(n5193), 
        .ZN(n5195) );
  ND4D1BWP U6641 ( .A1(n5192), .A2(n5191), .A3(n5190), .A4(n5189), .ZN(n5193)
         );
  AOI22D1BWP U6642 ( .A1(vectorData2[58]), .A2(n5188), .B1(vectorData2[234]), 
        .B2(n5187), .ZN(n5189) );
  AOI22D1BWP U6643 ( .A1(vectorData2[106]), .A2(n3671), .B1(vectorData2[74]), 
        .B2(n5186), .ZN(n5190) );
  AOI22D1BWP U6644 ( .A1(vectorData2[202]), .A2(n5227), .B1(vectorData2[42]), 
        .B2(n3601), .ZN(n5191) );
  AOI22D1BWP U6645 ( .A1(vectorData2[186]), .A2(n5233), .B1(vectorData2[138]), 
        .B2(n5226), .ZN(n5192) );
  AO22D1BWP U6646 ( .A1(vectorData2[154]), .A2(n5232), .B1(vectorData2[170]), 
        .B2(n5230), .Z(n5194) );
  AOI22D1BWP U6647 ( .A1(vectorData2[90]), .A2(n5185), .B1(vectorData2[250]), 
        .B2(n5229), .ZN(n5196) );
  AO222D1BWP U6648 ( .A1(n4550), .A2(n5501), .B1(n3650), .B2(n5408), .C1(
        vectorToLoad[93]), .C2(n4631), .Z(N4310) );
  NR2XD0BWP U6649 ( .A1(n5290), .A2(\intadd_34/A[2] ), .ZN(n5501) );
  AO222D1BWP U6650 ( .A1(n4550), .A2(n5504), .B1(n3650), .B2(n5410), .C1(
        vectorToLoad[94]), .C2(n3669), .Z(N4311) );
  NR2XD0BWP U6651 ( .A1(n5290), .A2(\intadd_34/A[3] ), .ZN(n5504) );
  AO222D1BWP U6652 ( .A1(n4550), .A2(n5507), .B1(n3650), .B2(n5412), .C1(
        vectorToLoad[95]), .C2(n3668), .Z(N4312) );
  NR2XD0BWP U6653 ( .A1(n5290), .A2(n6037), .ZN(n5507) );
  AO222D1BWP U6654 ( .A1(n3668), .A2(vectorToLoad[58]), .B1(n5403), .B2(n3649), 
        .C1(n4549), .C2(n5548), .Z(N4275) );
  AO222D1BWP U6655 ( .A1(n3669), .A2(vectorToLoad[96]), .B1(n3667), .B2(n5511), 
        .C1(n4548), .C2(n5512), .Z(N4313) );
  NR2XD0BWP U6656 ( .A1(n5370), .A2(n5813), .ZN(n5512) );
  AO211D1BWP U6657 ( .A1(instrIn[3]), .A2(n3928), .B(n3822), .C(n3821), .Z(
        N4195) );
  ND4D1BWP U6658 ( .A1(n3820), .A2(n3819), .A3(n3818), .A4(n3817), .ZN(n3821)
         );
  AOI22D1BWP U6659 ( .A1(n4687), .A2(vectorData2[35]), .B1(n4686), .B2(
        vectorData2[51]), .ZN(n3817) );
  AOI22D1BWP U6660 ( .A1(n4683), .A2(vectorData2[99]), .B1(n4685), .B2(
        vectorData2[19]), .ZN(n3818) );
  AOI22D1BWP U6661 ( .A1(n4682), .A2(vectorData2[67]), .B1(n4684), .B2(
        vectorData2[83]), .ZN(n3819) );
  AOI22D1BWP U6662 ( .A1(vectorData2[243]), .A2(n5229), .B1(vectorData2[115]), 
        .B2(n5231), .ZN(n5152) );
  AOI22D1BWP U6663 ( .A1(vectorData2[147]), .A2(n5232), .B1(vectorData2[211]), 
        .B2(n5228), .ZN(n5153) );
  AOI22D1BWP U6664 ( .A1(vectorData2[163]), .A2(n5230), .B1(vectorData2[179]), 
        .B2(n5233), .ZN(n5154) );
  AOI22D1BWP U6665 ( .A1(vectorData2[195]), .A2(n5227), .B1(vectorData2[131]), 
        .B2(n5226), .ZN(n5155) );
  AO22D1BWP U6666 ( .A1(n4681), .A2(vectorData2[3]), .B1(n4688), .B2(
        scalarData2[3]), .Z(n3822) );
  AO222D1BWP U6667 ( .A1(n3668), .A2(vectorToLoad[97]), .B1(n5515), .B2(n4628), 
        .C1(n3654), .C2(n5301), .Z(N4314) );
  AO222D1BWP U6668 ( .A1(n3669), .A2(vectorToLoad[57]), .B1(n5352), .B2(n3649), 
        .C1(n4549), .C2(n5547), .Z(N4274) );
  AO222D1BWP U6669 ( .A1(n3668), .A2(vectorToLoad[98]), .B1(n3654), .B2(n5304), 
        .C1(n5518), .C2(n4628), .Z(N4315) );
  AO222D1BWP U6670 ( .A1(n3669), .A2(vectorToLoad[99]), .B1(n3654), .B2(n5306), 
        .C1(n5521), .C2(n4628), .Z(N4316) );
  NR2XD0BWP U6671 ( .A1(n5292), .A2(n5291), .ZN(n5514) );
  AO211D1BWP U6672 ( .A1(instrIn[2]), .A2(n3928), .B(n5151), .C(n3807), .Z(
        N4194) );
  AOI31D1BWP U6673 ( .A1(n5144), .A2(n5146), .A3(n5145), .B(n3661), .ZN(n3807)
         );
  AOI22D1BWP U6674 ( .A1(vectorData2[130]), .A2(n5226), .B1(vectorData2[242]), 
        .B2(n5229), .ZN(n5145) );
  AOI22D1BWP U6675 ( .A1(vectorData2[146]), .A2(n5232), .B1(vectorData2[162]), 
        .B2(n5230), .ZN(n5146) );
  OA211D1BWP U6676 ( .A1(n5143), .A2(n3674), .B(n5142), .C(n5141), .Z(n5144)
         );
  AOI22D1BWP U6677 ( .A1(vectorData2[194]), .A2(n5227), .B1(vectorData2[178]), 
        .B2(n5233), .ZN(n5141) );
  AOI22D1BWP U6678 ( .A1(vectorData2[98]), .A2(n3671), .B1(vectorData2[210]), 
        .B2(n5228), .ZN(n5142) );
  ND4D1BWP U6679 ( .A1(n5150), .A2(n5149), .A3(n5148), .A4(n5147), .ZN(n5151)
         );
  AOI22D1BWP U6680 ( .A1(vectorData2[18]), .A2(n4685), .B1(scalarData2[2]), 
        .B2(n4688), .ZN(n5147) );
  AOI22D1BWP U6681 ( .A1(vectorData2[66]), .A2(n4682), .B1(vectorData2[34]), 
        .B2(n4687), .ZN(n5148) );
  AOI22D1BWP U6682 ( .A1(vectorData2[226]), .A2(n4694), .B1(vectorData2[2]), 
        .B2(n4681), .ZN(n5149) );
  AOI22D1BWP U6683 ( .A1(vectorData2[50]), .A2(n4686), .B1(vectorData2[82]), 
        .B2(n4684), .ZN(n5150) );
  OA211D1BWP U6684 ( .A1(n5299), .A2(n5509), .B(n5300), .C(n4403), .Z(n4404)
         );
  ND4D1BWP U6685 ( .A1(n5414), .A2(n4408), .A3(cycles[2]), .A4(n4402), .ZN(
        n4403) );
  AOI22D1BWP U6686 ( .A1(n3669), .A2(vectorToLoad[128]), .B1(n5297), .B2(n4626), .ZN(n5300) );
  OAI22D1BWP U6687 ( .A1(n4064), .A2(n3806), .B1(n3614), .B2(n3785), .ZN(N4134) );
  XNR2D1BWP U6688 ( .A1(n6004), .A2(n3679), .ZN(n3785) );
  AO222D1BWP U6689 ( .A1(n3668), .A2(vectorToLoad[56]), .B1(n5400), .B2(n3649), 
        .C1(n4549), .C2(n5546), .Z(N4273) );
  OAI211D1BWP U6690 ( .A1(n5517), .A2(n4405), .B(n5303), .C(n4535), .ZN(N4347)
         );
  AOI22D1BWP U6691 ( .A1(result[1]), .A2(n5331), .B1(n3668), .B2(
        vectorToLoad[129]), .ZN(n5303) );
  AO211D1BWP U6692 ( .A1(instrIn[1]), .A2(n3928), .B(n5140), .C(n3927), .Z(
        N4193) );
  AOI31D1BWP U6693 ( .A1(n5133), .A2(n5135), .A3(n5134), .B(n3661), .ZN(n3927)
         );
  AOI22D1BWP U6694 ( .A1(vectorData2[193]), .A2(n5227), .B1(vectorData2[113]), 
        .B2(n5231), .ZN(n5134) );
  AOI22D1BWP U6695 ( .A1(vectorData2[209]), .A2(n5228), .B1(vectorData2[241]), 
        .B2(n5229), .ZN(n5135) );
  OA211D1BWP U6696 ( .A1(n5132), .A2(n3673), .B(n5131), .C(n5130), .Z(n5133)
         );
  AOI22D1BWP U6697 ( .A1(vectorData2[145]), .A2(n5232), .B1(vectorData2[161]), 
        .B2(n5230), .ZN(n5130) );
  AOI22D1BWP U6698 ( .A1(vectorData2[33]), .A2(n3601), .B1(vectorData2[177]), 
        .B2(n5233), .ZN(n5131) );
  ND4D1BWP U6699 ( .A1(n5139), .A2(n5138), .A3(n5137), .A4(n5136), .ZN(n5140)
         );
  AOI22D1BWP U6700 ( .A1(vectorData2[17]), .A2(n4685), .B1(vectorData2[49]), 
        .B2(n4686), .ZN(n5136) );
  AOI22D1BWP U6701 ( .A1(vectorData2[225]), .A2(n4694), .B1(vectorData2[65]), 
        .B2(n4682), .ZN(n5137) );
  AOI22D1BWP U6702 ( .A1(vectorData2[1]), .A2(n4681), .B1(vectorData2[81]), 
        .B2(n4684), .ZN(n5138) );
  AOI22D1BWP U6703 ( .A1(vectorData2[97]), .A2(n4683), .B1(scalarData2[1]), 
        .B2(n4688), .ZN(n5139) );
  OAI211D1BWP U6704 ( .A1(n5520), .A2(n4405), .B(n5305), .C(n4535), .ZN(N4348)
         );
  AOI22D1BWP U6705 ( .A1(result[2]), .A2(n5331), .B1(n3668), .B2(
        vectorToLoad[130]), .ZN(n5305) );
  OAI211D1BWP U6706 ( .A1(n5523), .A2(n4405), .B(n5307), .C(n4535), .ZN(N4349)
         );
  AOI22D1BWP U6707 ( .A1(result[3]), .A2(n5331), .B1(n3668), .B2(
        vectorToLoad[131]), .ZN(n5307) );
  AO211D1BWP U6708 ( .A1(instrIn[0]), .A2(n3928), .B(n3758), .C(n3757), .Z(
        N4192) );
  ND4D1BWP U6709 ( .A1(n3756), .A2(n3755), .A3(n3754), .A4(n3753), .ZN(n3757)
         );
  AOI22D1BWP U6710 ( .A1(n4687), .A2(vectorData2[32]), .B1(n4686), .B2(
        vectorData2[48]), .ZN(n3753) );
  AOI22D1BWP U6711 ( .A1(n4683), .A2(vectorData2[96]), .B1(n4685), .B2(
        vectorData2[16]), .ZN(n3754) );
  AOI22D1BWP U6712 ( .A1(n4682), .A2(vectorData2[64]), .B1(n4684), .B2(
        vectorData2[80]), .ZN(n3755) );
  AOI22D1BWP U6713 ( .A1(vectorData2[176]), .A2(n5233), .B1(vectorData2[112]), 
        .B2(n5231), .ZN(n5125) );
  AOI22D1BWP U6714 ( .A1(vectorData2[160]), .A2(n5230), .B1(vectorData2[192]), 
        .B2(n5227), .ZN(n5126) );
  AOI22D1BWP U6715 ( .A1(vectorData2[128]), .A2(n5226), .B1(vectorData2[144]), 
        .B2(n5232), .ZN(n5127) );
  AOI22D1BWP U6716 ( .A1(vectorData2[208]), .A2(n5228), .B1(vectorData2[240]), 
        .B2(n5229), .ZN(n5128) );
  AO22D1BWP U6717 ( .A1(vectorData2[0]), .A2(n4681), .B1(scalarData2[0]), .B2(
        n4688), .Z(n3758) );
  OAI211D1BWP U6718 ( .A1(n5428), .A2(n4405), .B(n5309), .C(n4535), .ZN(N4350)
         );
  AOI22D1BWP U6719 ( .A1(result[4]), .A2(n5331), .B1(n3668), .B2(
        vectorToLoad[132]), .ZN(n5309) );
  AO222D1BWP U6720 ( .A1(n3668), .A2(vectorToLoad[55]), .B1(n5398), .B2(n3649), 
        .C1(n4549), .C2(n5545), .Z(N4272) );
  OAI211D1BWP U6721 ( .A1(n5431), .A2(n4405), .B(n5311), .C(n4535), .ZN(N4351)
         );
  AOI22D1BWP U6722 ( .A1(result[5]), .A2(n5331), .B1(n3668), .B2(
        vectorToLoad[133]), .ZN(n5311) );
  AO211D1BWP U6723 ( .A1(n4073), .A2(scalarData1[15]), .B(n3941), .C(n3940), 
        .Z(N4191) );
  AO22D1BWP U6724 ( .A1(n4072), .A2(vectorData1[15]), .B1(n4071), .B2(Addr[15]), .Z(n3940) );
  ND4D1BWP U6725 ( .A1(n7163), .A2(n7164), .A3(n7165), .A4(n7166), .ZN(
        vectorData1[15]) );
  AOI22D1BWP U6726 ( .A1(n3576), .A2(\vrf/regTable[5][15] ), .B1(n3567), .B2(
        \vrf/regTable[7][15] ), .ZN(n7166) );
  AOI22D1BWP U6727 ( .A1(n8285), .A2(\vrf/regTable[4][15] ), .B1(n3570), .B2(
        \vrf/regTable[6][15] ), .ZN(n7165) );
  AOI22D1BWP U6728 ( .A1(n3579), .A2(\vrf/regTable[1][15] ), .B1(n3575), .B2(
        \vrf/regTable[3][15] ), .ZN(n7164) );
  AOI22D1BWP U6729 ( .A1(n8278), .A2(\vrf/regTable[0][15] ), .B1(n3572), .B2(
        \vrf/regTable[2][15] ), .ZN(n7163) );
  AOI31D1BWP U6730 ( .A1(n5123), .A2(n5122), .A3(n5124), .B(n4070), .ZN(n3941)
         );
  AOI22D1BWP U6731 ( .A1(n5229), .A2(vectorData1[255]), .B1(n5232), .B2(
        vectorData1[159]), .ZN(n5124) );
  ND4D1BWP U6732 ( .A1(n7739), .A2(n7740), .A3(n7741), .A4(n7742), .ZN(
        vectorData1[159]) );
  AOI22D1BWP U6733 ( .A1(n3576), .A2(\vrf/regTable[5][159] ), .B1(n3595), .B2(
        \vrf/regTable[7][159] ), .ZN(n7742) );
  AOI22D1BWP U6734 ( .A1(n3574), .A2(\vrf/regTable[4][159] ), .B1(n3596), .B2(
        \vrf/regTable[6][159] ), .ZN(n7741) );
  AOI22D1BWP U6735 ( .A1(n3579), .A2(\vrf/regTable[1][159] ), .B1(n3575), .B2(
        \vrf/regTable[3][159] ), .ZN(n7740) );
  AOI22D1BWP U6736 ( .A1(n3581), .A2(\vrf/regTable[0][159] ), .B1(n3594), .B2(
        \vrf/regTable[2][159] ), .ZN(n7739) );
  ND4D1BWP U6737 ( .A1(n8123), .A2(n8124), .A3(n8125), .A4(n8126), .ZN(
        vectorData1[255]) );
  AOI22D1BWP U6738 ( .A1(n3576), .A2(\vrf/regTable[5][255] ), .B1(n3567), .B2(
        \vrf/regTable[7][255] ), .ZN(n8126) );
  AOI22D1BWP U6739 ( .A1(n3574), .A2(\vrf/regTable[4][255] ), .B1(n3570), .B2(
        \vrf/regTable[6][255] ), .ZN(n8125) );
  AOI22D1BWP U6740 ( .A1(n3579), .A2(\vrf/regTable[1][255] ), .B1(n3575), .B2(
        \vrf/regTable[3][255] ), .ZN(n8124) );
  AOI22D1BWP U6741 ( .A1(n3581), .A2(\vrf/regTable[0][255] ), .B1(n3572), .B2(
        \vrf/regTable[2][255] ), .ZN(n8123) );
  AOI211XD0BWP U6742 ( .A1(n5226), .A2(vectorData1[143]), .B(n5121), .C(n5120), 
        .ZN(n5122) );
  ND4D1BWP U6743 ( .A1(n5119), .A2(n5118), .A3(n5117), .A4(n5116), .ZN(n5120)
         );
  AOI22D1BWP U6744 ( .A1(n3601), .A2(vectorData1[47]), .B1(n5188), .B2(
        vectorData1[63]), .ZN(n5116) );
  ND4D1BWP U6745 ( .A1(n7355), .A2(n7356), .A3(n7357), .A4(n7358), .ZN(
        vectorData1[63]) );
  AOI22D1BWP U6746 ( .A1(n3576), .A2(\vrf/regTable[5][63] ), .B1(n3567), .B2(
        \vrf/regTable[7][63] ), .ZN(n7358) );
  AOI22D1BWP U6747 ( .A1(n3574), .A2(\vrf/regTable[4][63] ), .B1(n3570), .B2(
        \vrf/regTable[6][63] ), .ZN(n7357) );
  AOI22D1BWP U6748 ( .A1(n3579), .A2(\vrf/regTable[1][63] ), .B1(n3575), .B2(
        \vrf/regTable[3][63] ), .ZN(n7356) );
  AOI22D1BWP U6749 ( .A1(n3581), .A2(\vrf/regTable[0][63] ), .B1(n3572), .B2(
        \vrf/regTable[2][63] ), .ZN(n7355) );
  ND4D1BWP U6750 ( .A1(n7291), .A2(n7292), .A3(n7293), .A4(n7294), .ZN(
        vectorData1[47]) );
  AOI22D1BWP U6751 ( .A1(n3576), .A2(\vrf/regTable[5][47] ), .B1(n3595), .B2(
        \vrf/regTable[7][47] ), .ZN(n7294) );
  AOI22D1BWP U6752 ( .A1(n3574), .A2(\vrf/regTable[4][47] ), .B1(n3596), .B2(
        \vrf/regTable[6][47] ), .ZN(n7293) );
  AOI22D1BWP U6753 ( .A1(n3579), .A2(\vrf/regTable[1][47] ), .B1(n3599), .B2(
        \vrf/regTable[3][47] ), .ZN(n7292) );
  AOI22D1BWP U6754 ( .A1(n3581), .A2(\vrf/regTable[0][47] ), .B1(n3594), .B2(
        \vrf/regTable[2][47] ), .ZN(n7291) );
  AOI22D1BWP U6755 ( .A1(n5185), .A2(vectorData1[95]), .B1(n5184), .B2(
        vectorData1[31]), .ZN(n5117) );
  ND4D1BWP U6756 ( .A1(n7227), .A2(n7228), .A3(n7229), .A4(n7230), .ZN(
        vectorData1[31]) );
  AOI22D1BWP U6757 ( .A1(n3576), .A2(\vrf/regTable[5][31] ), .B1(n3567), .B2(
        \vrf/regTable[7][31] ), .ZN(n7230) );
  AOI22D1BWP U6758 ( .A1(n3574), .A2(\vrf/regTable[4][31] ), .B1(n3570), .B2(
        \vrf/regTable[6][31] ), .ZN(n7229) );
  AOI22D1BWP U6759 ( .A1(n3579), .A2(\vrf/regTable[1][31] ), .B1(n3575), .B2(
        \vrf/regTable[3][31] ), .ZN(n7228) );
  AOI22D1BWP U6760 ( .A1(n3581), .A2(\vrf/regTable[0][31] ), .B1(n3572), .B2(
        \vrf/regTable[2][31] ), .ZN(n7227) );
  ND4D1BWP U6761 ( .A1(n7483), .A2(n7484), .A3(n7485), .A4(n7486), .ZN(
        vectorData1[95]) );
  AOI22D1BWP U6762 ( .A1(n3576), .A2(\vrf/regTable[5][95] ), .B1(n3567), .B2(
        \vrf/regTable[7][95] ), .ZN(n7486) );
  AOI22D1BWP U6763 ( .A1(n3574), .A2(\vrf/regTable[4][95] ), .B1(n3570), .B2(
        \vrf/regTable[6][95] ), .ZN(n7485) );
  AOI22D1BWP U6764 ( .A1(n3579), .A2(\vrf/regTable[1][95] ), .B1(n3575), .B2(
        \vrf/regTable[3][95] ), .ZN(n7484) );
  AOI22D1BWP U6765 ( .A1(n3581), .A2(\vrf/regTable[0][95] ), .B1(n3572), .B2(
        \vrf/regTable[2][95] ), .ZN(n7483) );
  AOI22D1BWP U6766 ( .A1(n5230), .A2(vectorData1[175]), .B1(n5227), .B2(
        vectorData1[207]), .ZN(n5118) );
  ND4D1BWP U6767 ( .A1(n7931), .A2(n7932), .A3(n7933), .A4(n7934), .ZN(
        vectorData1[207]) );
  AOI22D1BWP U6768 ( .A1(n3576), .A2(\vrf/regTable[5][207] ), .B1(n3595), .B2(
        \vrf/regTable[7][207] ), .ZN(n7934) );
  AOI22D1BWP U6769 ( .A1(n3574), .A2(\vrf/regTable[4][207] ), .B1(n3596), .B2(
        \vrf/regTable[6][207] ), .ZN(n7933) );
  AOI22D1BWP U6770 ( .A1(n3579), .A2(\vrf/regTable[1][207] ), .B1(n3599), .B2(
        \vrf/regTable[3][207] ), .ZN(n7932) );
  AOI22D1BWP U6771 ( .A1(n3581), .A2(\vrf/regTable[0][207] ), .B1(n3594), .B2(
        \vrf/regTable[2][207] ), .ZN(n7931) );
  ND4D1BWP U6772 ( .A1(n7803), .A2(n7804), .A3(n7805), .A4(n7806), .ZN(
        vectorData1[175]) );
  AOI22D1BWP U6773 ( .A1(n3576), .A2(\vrf/regTable[5][175] ), .B1(n3567), .B2(
        \vrf/regTable[7][175] ), .ZN(n7806) );
  AOI22D1BWP U6774 ( .A1(n3574), .A2(\vrf/regTable[4][175] ), .B1(n3570), .B2(
        \vrf/regTable[6][175] ), .ZN(n7805) );
  AOI22D1BWP U6775 ( .A1(n3579), .A2(\vrf/regTable[1][175] ), .B1(n3575), .B2(
        \vrf/regTable[3][175] ), .ZN(n7804) );
  AOI22D1BWP U6776 ( .A1(n3581), .A2(\vrf/regTable[0][175] ), .B1(n3572), .B2(
        \vrf/regTable[2][175] ), .ZN(n7803) );
  AOI22D1BWP U6777 ( .A1(n5187), .A2(vectorData1[239]), .B1(n5231), .B2(
        vectorData1[127]), .ZN(n5119) );
  ND4D1BWP U6778 ( .A1(n7611), .A2(n7612), .A3(n7613), .A4(n7614), .ZN(
        vectorData1[127]) );
  AOI22D1BWP U6779 ( .A1(n3576), .A2(\vrf/regTable[5][127] ), .B1(n3567), .B2(
        \vrf/regTable[7][127] ), .ZN(n7614) );
  AOI22D1BWP U6780 ( .A1(n3574), .A2(\vrf/regTable[4][127] ), .B1(n3570), .B2(
        \vrf/regTable[6][127] ), .ZN(n7613) );
  AOI22D1BWP U6781 ( .A1(n3579), .A2(\vrf/regTable[1][127] ), .B1(n3599), .B2(
        \vrf/regTable[3][127] ), .ZN(n7612) );
  AOI22D1BWP U6782 ( .A1(n3581), .A2(\vrf/regTable[0][127] ), .B1(n3572), .B2(
        \vrf/regTable[2][127] ), .ZN(n7611) );
  ND4D1BWP U6783 ( .A1(n8059), .A2(n8060), .A3(n8061), .A4(n8062), .ZN(
        vectorData1[239]) );
  AOI22D1BWP U6784 ( .A1(n3576), .A2(\vrf/regTable[5][239] ), .B1(n3595), .B2(
        \vrf/regTable[7][239] ), .ZN(n8062) );
  AOI22D1BWP U6785 ( .A1(n8285), .A2(\vrf/regTable[4][239] ), .B1(n3596), .B2(
        \vrf/regTable[6][239] ), .ZN(n8061) );
  AOI22D1BWP U6786 ( .A1(n3579), .A2(\vrf/regTable[1][239] ), .B1(n3599), .B2(
        \vrf/regTable[3][239] ), .ZN(n8060) );
  AOI22D1BWP U6787 ( .A1(n8278), .A2(\vrf/regTable[0][239] ), .B1(n3594), .B2(
        \vrf/regTable[2][239] ), .ZN(n8059) );
  AO22D1BWP U6788 ( .A1(n3671), .A2(vectorData1[111]), .B1(n5186), .B2(
        vectorData1[79]), .Z(n5121) );
  ND4D1BWP U6789 ( .A1(n7419), .A2(n7420), .A3(n7421), .A4(n7422), .ZN(
        vectorData1[79]) );
  AOI22D1BWP U6790 ( .A1(n3576), .A2(\vrf/regTable[5][79] ), .B1(n3567), .B2(
        \vrf/regTable[7][79] ), .ZN(n7422) );
  AOI22D1BWP U6791 ( .A1(n7115), .A2(\vrf/regTable[4][79] ), .B1(n3570), .B2(
        \vrf/regTable[6][79] ), .ZN(n7421) );
  AOI22D1BWP U6792 ( .A1(n3579), .A2(\vrf/regTable[1][79] ), .B1(n3575), .B2(
        \vrf/regTable[3][79] ), .ZN(n7420) );
  AOI22D1BWP U6793 ( .A1(n7108), .A2(\vrf/regTable[0][79] ), .B1(n3572), .B2(
        \vrf/regTable[2][79] ), .ZN(n7419) );
  ND4D1BWP U6794 ( .A1(n7547), .A2(n7548), .A3(n7549), .A4(n7550), .ZN(
        vectorData1[111]) );
  AOI22D1BWP U6795 ( .A1(n3576), .A2(\vrf/regTable[5][111] ), .B1(n3595), .B2(
        \vrf/regTable[7][111] ), .ZN(n7550) );
  AOI22D1BWP U6796 ( .A1(n7115), .A2(\vrf/regTable[4][111] ), .B1(n3596), .B2(
        \vrf/regTable[6][111] ), .ZN(n7549) );
  AOI22D1BWP U6797 ( .A1(n3579), .A2(\vrf/regTable[1][111] ), .B1(n3599), .B2(
        \vrf/regTable[3][111] ), .ZN(n7548) );
  AOI22D1BWP U6798 ( .A1(n7108), .A2(\vrf/regTable[0][111] ), .B1(n3594), .B2(
        \vrf/regTable[2][111] ), .ZN(n7547) );
  ND4D1BWP U6799 ( .A1(n7675), .A2(n7676), .A3(n7677), .A4(n7678), .ZN(
        vectorData1[143]) );
  AOI22D1BWP U6800 ( .A1(n3576), .A2(\vrf/regTable[5][143] ), .B1(n3567), .B2(
        \vrf/regTable[7][143] ), .ZN(n7678) );
  AOI22D1BWP U6801 ( .A1(n3574), .A2(\vrf/regTable[4][143] ), .B1(n3570), .B2(
        \vrf/regTable[6][143] ), .ZN(n7677) );
  AOI22D1BWP U6802 ( .A1(n3579), .A2(\vrf/regTable[1][143] ), .B1(n3599), .B2(
        \vrf/regTable[3][143] ), .ZN(n7676) );
  AOI22D1BWP U6803 ( .A1(n3581), .A2(\vrf/regTable[0][143] ), .B1(n3572), .B2(
        \vrf/regTable[2][143] ), .ZN(n7675) );
  AOI22D1BWP U6804 ( .A1(n5228), .A2(vectorData1[223]), .B1(n5233), .B2(
        vectorData1[191]), .ZN(n5123) );
  ND4D1BWP U6805 ( .A1(n7867), .A2(n7868), .A3(n7869), .A4(n7870), .ZN(
        vectorData1[191]) );
  AOI22D1BWP U6806 ( .A1(n3576), .A2(\vrf/regTable[5][191] ), .B1(n3595), .B2(
        \vrf/regTable[7][191] ), .ZN(n7870) );
  AOI22D1BWP U6807 ( .A1(n3574), .A2(\vrf/regTable[4][191] ), .B1(n3596), .B2(
        \vrf/regTable[6][191] ), .ZN(n7869) );
  AOI22D1BWP U6808 ( .A1(n3579), .A2(\vrf/regTable[1][191] ), .B1(n3599), .B2(
        \vrf/regTable[3][191] ), .ZN(n7868) );
  AOI22D1BWP U6809 ( .A1(n3581), .A2(\vrf/regTable[0][191] ), .B1(n3594), .B2(
        \vrf/regTable[2][191] ), .ZN(n7867) );
  ND4D1BWP U6810 ( .A1(n7995), .A2(n7996), .A3(n7997), .A4(n7998), .ZN(
        vectorData1[223]) );
  AOI22D1BWP U6811 ( .A1(n3576), .A2(\vrf/regTable[5][223] ), .B1(n3567), .B2(
        \vrf/regTable[7][223] ), .ZN(n7998) );
  AOI22D1BWP U6812 ( .A1(n8285), .A2(\vrf/regTable[4][223] ), .B1(n3570), .B2(
        \vrf/regTable[6][223] ), .ZN(n7997) );
  AOI22D1BWP U6813 ( .A1(n3579), .A2(\vrf/regTable[1][223] ), .B1(n3575), .B2(
        \vrf/regTable[3][223] ), .ZN(n7996) );
  AOI22D1BWP U6814 ( .A1(n8278), .A2(\vrf/regTable[0][223] ), .B1(n3572), .B2(
        \vrf/regTable[2][223] ), .ZN(n7995) );
  ND4D1BWP U6815 ( .A1(n8333), .A2(n8334), .A3(n8335), .A4(n8336), .ZN(
        scalarData1[15]) );
  AOI22D1BWP U6816 ( .A1(n8287), .A2(\srf/regTable[5][15] ), .B1(n8288), .B2(
        \srf/regTable[7][15] ), .ZN(n8336) );
  AOI22D1BWP U6817 ( .A1(n8285), .A2(\srf/regTable[4][15] ), .B1(n8286), .B2(
        \srf/regTable[6][15] ), .ZN(n8335) );
  AOI22D1BWP U6818 ( .A1(n8282), .A2(\srf/regTable[1][15] ), .B1(n8284), .B2(
        \srf/regTable[3][15] ), .ZN(n8334) );
  AOI22D1BWP U6819 ( .A1(n8278), .A2(\srf/regTable[0][15] ), .B1(n8280), .B2(
        \srf/regTable[2][15] ), .ZN(n8333) );
  OAI211D1BWP U6820 ( .A1(n5434), .A2(n4405), .B(n5313), .C(n4535), .ZN(N4352)
         );
  AOI22D1BWP U6821 ( .A1(result[6]), .A2(n5331), .B1(n3668), .B2(
        vectorToLoad[134]), .ZN(n5313) );
  AO222D1BWP U6822 ( .A1(n3635), .A2(n4548), .B1(n5524), .B2(n3667), .C1(n3669), .C2(vectorToLoad[100]), .Z(N4317) );
  AO222D1BWP U6823 ( .A1(n3669), .A2(vectorToLoad[54]), .B1(n5396), .B2(n3649), 
        .C1(n4549), .C2(n5544), .Z(N4271) );
  OAI211D1BWP U6824 ( .A1(n5437), .A2(n4405), .B(n5315), .C(n4535), .ZN(N4353)
         );
  AOI22D1BWP U6825 ( .A1(result[7]), .A2(n5331), .B1(n3668), .B2(
        vectorToLoad[135]), .ZN(n5315) );
  ND4D1BWP U6826 ( .A1(n7863), .A2(n7864), .A3(n7865), .A4(n7866), .ZN(
        vectorData1[190]) );
  AOI22D1BWP U6827 ( .A1(n3576), .A2(\vrf/regTable[5][190] ), .B1(n3595), .B2(
        \vrf/regTable[7][190] ), .ZN(n7866) );
  AOI22D1BWP U6828 ( .A1(n3574), .A2(\vrf/regTable[4][190] ), .B1(n3596), .B2(
        \vrf/regTable[6][190] ), .ZN(n7865) );
  AOI22D1BWP U6829 ( .A1(n3579), .A2(\vrf/regTable[1][190] ), .B1(n3599), .B2(
        \vrf/regTable[3][190] ), .ZN(n7864) );
  AOI22D1BWP U6830 ( .A1(n3581), .A2(\vrf/regTable[0][190] ), .B1(n3594), .B2(
        \vrf/regTable[2][190] ), .ZN(n7863) );
  AOI22D1BWP U6831 ( .A1(n3576), .A2(\vrf/regTable[5][238] ), .B1(n3595), .B2(
        \vrf/regTable[7][238] ), .ZN(n8058) );
  AOI22D1BWP U6832 ( .A1(n7115), .A2(\vrf/regTable[4][238] ), .B1(n3596), .B2(
        \vrf/regTable[6][238] ), .ZN(n8057) );
  AOI22D1BWP U6833 ( .A1(n3579), .A2(\vrf/regTable[1][238] ), .B1(n3599), .B2(
        \vrf/regTable[3][238] ), .ZN(n8056) );
  AOI22D1BWP U6834 ( .A1(n7108), .A2(\vrf/regTable[0][238] ), .B1(n3594), .B2(
        \vrf/regTable[2][238] ), .ZN(n8055) );
  AOI22D1BWP U6835 ( .A1(n5226), .A2(vectorData1[142]), .B1(n5227), .B2(
        vectorData1[206]), .ZN(n5112) );
  ND4D1BWP U6836 ( .A1(n7927), .A2(n7928), .A3(n7929), .A4(n7930), .ZN(
        vectorData1[206]) );
  AOI22D1BWP U6837 ( .A1(n3576), .A2(\vrf/regTable[5][206] ), .B1(n3567), .B2(
        \vrf/regTable[7][206] ), .ZN(n7930) );
  AOI22D1BWP U6838 ( .A1(n3574), .A2(\vrf/regTable[4][206] ), .B1(n3570), .B2(
        \vrf/regTable[6][206] ), .ZN(n7929) );
  AOI22D1BWP U6839 ( .A1(n3579), .A2(\vrf/regTable[1][206] ), .B1(n3575), .B2(
        \vrf/regTable[3][206] ), .ZN(n7928) );
  AOI22D1BWP U6840 ( .A1(n3581), .A2(\vrf/regTable[0][206] ), .B1(n3572), .B2(
        \vrf/regTable[2][206] ), .ZN(n7927) );
  ND4D1BWP U6841 ( .A1(n7671), .A2(n7672), .A3(n7673), .A4(n7674), .ZN(
        vectorData1[142]) );
  AOI22D1BWP U6842 ( .A1(n3576), .A2(\vrf/regTable[5][142] ), .B1(n3595), .B2(
        \vrf/regTable[7][142] ), .ZN(n7674) );
  AOI22D1BWP U6843 ( .A1(n3574), .A2(\vrf/regTable[4][142] ), .B1(n3596), .B2(
        \vrf/regTable[6][142] ), .ZN(n7673) );
  AOI22D1BWP U6844 ( .A1(n3579), .A2(\vrf/regTable[1][142] ), .B1(n3599), .B2(
        \vrf/regTable[3][142] ), .ZN(n7672) );
  AOI22D1BWP U6845 ( .A1(n3581), .A2(\vrf/regTable[0][142] ), .B1(n3594), .B2(
        \vrf/regTable[2][142] ), .ZN(n7671) );
  AOI22D1BWP U6846 ( .A1(n5231), .A2(vectorData1[126]), .B1(n5184), .B2(
        vectorData1[30]), .ZN(n5113) );
  ND4D1BWP U6847 ( .A1(n7223), .A2(n7224), .A3(n7225), .A4(n7226), .ZN(
        vectorData1[30]) );
  AOI22D1BWP U6848 ( .A1(n3576), .A2(\vrf/regTable[5][30] ), .B1(n3567), .B2(
        \vrf/regTable[7][30] ), .ZN(n7226) );
  AOI22D1BWP U6849 ( .A1(n8285), .A2(\vrf/regTable[4][30] ), .B1(n3570), .B2(
        \vrf/regTable[6][30] ), .ZN(n7225) );
  AOI22D1BWP U6850 ( .A1(n3579), .A2(\vrf/regTable[1][30] ), .B1(n3575), .B2(
        \vrf/regTable[3][30] ), .ZN(n7224) );
  AOI22D1BWP U6851 ( .A1(n8278), .A2(\vrf/regTable[0][30] ), .B1(n3572), .B2(
        \vrf/regTable[2][30] ), .ZN(n7223) );
  ND4D1BWP U6852 ( .A1(n7607), .A2(n7608), .A3(n7609), .A4(n7610), .ZN(
        vectorData1[126]) );
  AOI22D1BWP U6853 ( .A1(n3576), .A2(\vrf/regTable[5][126] ), .B1(n3567), .B2(
        \vrf/regTable[7][126] ), .ZN(n7610) );
  AOI22D1BWP U6854 ( .A1(n3574), .A2(\vrf/regTable[4][126] ), .B1(n3570), .B2(
        \vrf/regTable[6][126] ), .ZN(n7609) );
  AOI22D1BWP U6855 ( .A1(n3579), .A2(\vrf/regTable[1][126] ), .B1(n3575), .B2(
        \vrf/regTable[3][126] ), .ZN(n7608) );
  AOI22D1BWP U6856 ( .A1(n3581), .A2(\vrf/regTable[0][126] ), .B1(n3572), .B2(
        \vrf/regTable[2][126] ), .ZN(n7607) );
  AOI22D1BWP U6857 ( .A1(n3671), .A2(vectorData1[110]), .B1(n3601), .B2(
        vectorData1[46]), .ZN(n5114) );
  ND4D1BWP U6858 ( .A1(n7287), .A2(n7288), .A3(n7289), .A4(n7290), .ZN(
        vectorData1[46]) );
  AOI22D1BWP U6859 ( .A1(n3576), .A2(\vrf/regTable[5][46] ), .B1(n3595), .B2(
        \vrf/regTable[7][46] ), .ZN(n7290) );
  AOI22D1BWP U6860 ( .A1(n3574), .A2(\vrf/regTable[4][46] ), .B1(n3596), .B2(
        \vrf/regTable[6][46] ), .ZN(n7289) );
  AOI22D1BWP U6861 ( .A1(n3579), .A2(\vrf/regTable[1][46] ), .B1(n3599), .B2(
        \vrf/regTable[3][46] ), .ZN(n7288) );
  AOI22D1BWP U6862 ( .A1(n3581), .A2(\vrf/regTable[0][46] ), .B1(n3594), .B2(
        \vrf/regTable[2][46] ), .ZN(n7287) );
  ND4D1BWP U6863 ( .A1(n7543), .A2(n7544), .A3(n7545), .A4(n7546), .ZN(
        vectorData1[110]) );
  AOI22D1BWP U6864 ( .A1(n3576), .A2(\vrf/regTable[5][110] ), .B1(n3595), .B2(
        \vrf/regTable[7][110] ), .ZN(n7546) );
  AOI22D1BWP U6865 ( .A1(n3574), .A2(\vrf/regTable[4][110] ), .B1(n3596), .B2(
        \vrf/regTable[6][110] ), .ZN(n7545) );
  AOI22D1BWP U6866 ( .A1(n3579), .A2(\vrf/regTable[1][110] ), .B1(n3599), .B2(
        \vrf/regTable[3][110] ), .ZN(n7544) );
  AOI22D1BWP U6867 ( .A1(n3581), .A2(\vrf/regTable[0][110] ), .B1(n3594), .B2(
        \vrf/regTable[2][110] ), .ZN(n7543) );
  AOI22D1BWP U6868 ( .A1(n5229), .A2(vectorData1[254]), .B1(n5188), .B2(
        vectorData1[62]), .ZN(n5115) );
  ND4D1BWP U6869 ( .A1(n7351), .A2(n7352), .A3(n7353), .A4(n7354), .ZN(
        vectorData1[62]) );
  AOI22D1BWP U6870 ( .A1(n3576), .A2(\vrf/regTable[5][62] ), .B1(n3567), .B2(
        \vrf/regTable[7][62] ), .ZN(n7354) );
  AOI22D1BWP U6871 ( .A1(n3574), .A2(\vrf/regTable[4][62] ), .B1(n3570), .B2(
        \vrf/regTable[6][62] ), .ZN(n7353) );
  AOI22D1BWP U6872 ( .A1(n3579), .A2(\vrf/regTable[1][62] ), .B1(n3575), .B2(
        \vrf/regTable[3][62] ), .ZN(n7352) );
  AOI22D1BWP U6873 ( .A1(n3581), .A2(\vrf/regTable[0][62] ), .B1(n3572), .B2(
        \vrf/regTable[2][62] ), .ZN(n7351) );
  ND4D1BWP U6874 ( .A1(n8119), .A2(n8120), .A3(n8121), .A4(n8122), .ZN(
        vectorData1[254]) );
  AOI22D1BWP U6875 ( .A1(n3576), .A2(\vrf/regTable[5][254] ), .B1(n7118), .B2(
        \vrf/regTable[7][254] ), .ZN(n8122) );
  AOI22D1BWP U6876 ( .A1(n3574), .A2(\vrf/regTable[4][254] ), .B1(n7116), .B2(
        \vrf/regTable[6][254] ), .ZN(n8121) );
  AOI22D1BWP U6877 ( .A1(n3579), .A2(\vrf/regTable[1][254] ), .B1(n7114), .B2(
        \vrf/regTable[3][254] ), .ZN(n8120) );
  AOI22D1BWP U6878 ( .A1(n3581), .A2(\vrf/regTable[0][254] ), .B1(n7110), .B2(
        \vrf/regTable[2][254] ), .ZN(n8119) );
  ND4D1BWP U6879 ( .A1(n7415), .A2(n7416), .A3(n7417), .A4(n7418), .ZN(
        vectorData1[78]) );
  AOI22D1BWP U6880 ( .A1(n7117), .A2(\vrf/regTable[5][78] ), .B1(n3595), .B2(
        \vrf/regTable[7][78] ), .ZN(n7418) );
  AOI22D1BWP U6881 ( .A1(n7115), .A2(\vrf/regTable[4][78] ), .B1(n3596), .B2(
        \vrf/regTable[6][78] ), .ZN(n7417) );
  AOI22D1BWP U6882 ( .A1(n7112), .A2(\vrf/regTable[1][78] ), .B1(n3599), .B2(
        \vrf/regTable[3][78] ), .ZN(n7416) );
  AOI22D1BWP U6883 ( .A1(n7108), .A2(\vrf/regTable[0][78] ), .B1(n3594), .B2(
        \vrf/regTable[2][78] ), .ZN(n7415) );
  ND4D1BWP U6884 ( .A1(n7799), .A2(n7800), .A3(n7801), .A4(n7802), .ZN(
        vectorData1[174]) );
  AOI22D1BWP U6885 ( .A1(n3576), .A2(\vrf/regTable[5][174] ), .B1(n3595), .B2(
        \vrf/regTable[7][174] ), .ZN(n7802) );
  AOI22D1BWP U6886 ( .A1(n3574), .A2(\vrf/regTable[4][174] ), .B1(n3596), .B2(
        \vrf/regTable[6][174] ), .ZN(n7801) );
  AOI22D1BWP U6887 ( .A1(n3579), .A2(\vrf/regTable[1][174] ), .B1(n3599), .B2(
        \vrf/regTable[3][174] ), .ZN(n7800) );
  AOI22D1BWP U6888 ( .A1(n3581), .A2(\vrf/regTable[0][174] ), .B1(n3594), .B2(
        \vrf/regTable[2][174] ), .ZN(n7799) );
  AOI22D1BWP U6889 ( .A1(n3576), .A2(\vrf/regTable[5][222] ), .B1(n3595), .B2(
        \vrf/regTable[7][222] ), .ZN(n7994) );
  AOI22D1BWP U6890 ( .A1(n3574), .A2(\vrf/regTable[4][222] ), .B1(n3596), .B2(
        \vrf/regTable[6][222] ), .ZN(n7993) );
  AOI22D1BWP U6891 ( .A1(n3579), .A2(\vrf/regTable[1][222] ), .B1(n3599), .B2(
        \vrf/regTable[3][222] ), .ZN(n7992) );
  AOI22D1BWP U6892 ( .A1(n3581), .A2(\vrf/regTable[0][222] ), .B1(n3594), .B2(
        \vrf/regTable[2][222] ), .ZN(n7991) );
  ND4D1BWP U6893 ( .A1(n7735), .A2(n7736), .A3(n7737), .A4(n7738), .ZN(
        vectorData1[158]) );
  AOI22D1BWP U6894 ( .A1(n3576), .A2(\vrf/regTable[5][158] ), .B1(n3567), .B2(
        \vrf/regTable[7][158] ), .ZN(n7738) );
  AOI22D1BWP U6895 ( .A1(n3574), .A2(\vrf/regTable[4][158] ), .B1(n3570), .B2(
        \vrf/regTable[6][158] ), .ZN(n7737) );
  AOI22D1BWP U6896 ( .A1(n3579), .A2(\vrf/regTable[1][158] ), .B1(n3599), .B2(
        \vrf/regTable[3][158] ), .ZN(n7736) );
  AOI22D1BWP U6897 ( .A1(n3581), .A2(\vrf/regTable[0][158] ), .B1(n3572), .B2(
        \vrf/regTable[2][158] ), .ZN(n7735) );
  ND4D1BWP U6898 ( .A1(n7479), .A2(n7480), .A3(n7481), .A4(n7482), .ZN(
        vectorData1[94]) );
  AOI22D1BWP U6899 ( .A1(n7117), .A2(\vrf/regTable[5][94] ), .B1(n3567), .B2(
        \vrf/regTable[7][94] ), .ZN(n7482) );
  AOI22D1BWP U6900 ( .A1(n7115), .A2(\vrf/regTable[4][94] ), .B1(n3570), .B2(
        \vrf/regTable[6][94] ), .ZN(n7481) );
  AOI22D1BWP U6901 ( .A1(n7112), .A2(\vrf/regTable[1][94] ), .B1(n3575), .B2(
        \vrf/regTable[3][94] ), .ZN(n7480) );
  AOI22D1BWP U6902 ( .A1(n7108), .A2(\vrf/regTable[0][94] ), .B1(n3572), .B2(
        \vrf/regTable[2][94] ), .ZN(n7479) );
  OAI211D1BWP U6903 ( .A1(n5440), .A2(n4405), .B(n5317), .C(n4535), .ZN(N4354)
         );
  AOI22D1BWP U6904 ( .A1(result[8]), .A2(n5331), .B1(n3668), .B2(
        vectorToLoad[136]), .ZN(n5317) );
  AO211D1BWP U6905 ( .A1(n4073), .A2(scalarData1[12]), .B(n3863), .C(n3862), 
        .Z(N4188) );
  AO22D1BWP U6906 ( .A1(n4072), .A2(vectorData1[12]), .B1(n4071), .B2(Addr[12]), .Z(n3862) );
  ND4D1BWP U6907 ( .A1(n7155), .A2(n7156), .A3(n7157), .A4(n7158), .ZN(
        vectorData1[12]) );
  AOI22D1BWP U6908 ( .A1(n3576), .A2(\vrf/regTable[5][12] ), .B1(n3595), .B2(
        \vrf/regTable[7][12] ), .ZN(n7158) );
  AOI22D1BWP U6909 ( .A1(n7115), .A2(\vrf/regTable[4][12] ), .B1(n3596), .B2(
        \vrf/regTable[6][12] ), .ZN(n7157) );
  AOI22D1BWP U6910 ( .A1(n3579), .A2(\vrf/regTable[1][12] ), .B1(n3599), .B2(
        \vrf/regTable[3][12] ), .ZN(n7156) );
  AOI22D1BWP U6911 ( .A1(n7108), .A2(\vrf/regTable[0][12] ), .B1(n3594), .B2(
        \vrf/regTable[2][12] ), .ZN(n7155) );
  AOI31D1BWP U6912 ( .A1(n5101), .A2(n5100), .A3(n5102), .B(n4070), .ZN(n3863)
         );
  AOI22D1BWP U6913 ( .A1(n5229), .A2(vectorData1[252]), .B1(n5230), .B2(
        vectorData1[172]), .ZN(n5102) );
  ND4D1BWP U6914 ( .A1(n7791), .A2(n7792), .A3(n7793), .A4(n7794), .ZN(
        vectorData1[172]) );
  AOI22D1BWP U6915 ( .A1(n3576), .A2(\vrf/regTable[5][172] ), .B1(n3595), .B2(
        \vrf/regTable[7][172] ), .ZN(n7794) );
  AOI22D1BWP U6916 ( .A1(n3574), .A2(\vrf/regTable[4][172] ), .B1(n3596), .B2(
        \vrf/regTable[6][172] ), .ZN(n7793) );
  AOI22D1BWP U6917 ( .A1(n3579), .A2(\vrf/regTable[1][172] ), .B1(n3599), .B2(
        \vrf/regTable[3][172] ), .ZN(n7792) );
  AOI22D1BWP U6918 ( .A1(n3581), .A2(\vrf/regTable[0][172] ), .B1(n3594), .B2(
        \vrf/regTable[2][172] ), .ZN(n7791) );
  ND4D1BWP U6919 ( .A1(n8111), .A2(n8112), .A3(n8113), .A4(n8114), .ZN(
        vectorData1[252]) );
  AOI22D1BWP U6920 ( .A1(n3576), .A2(\vrf/regTable[5][252] ), .B1(n7118), .B2(
        \vrf/regTable[7][252] ), .ZN(n8114) );
  AOI22D1BWP U6921 ( .A1(n8285), .A2(\vrf/regTable[4][252] ), .B1(n7116), .B2(
        \vrf/regTable[6][252] ), .ZN(n8113) );
  AOI22D1BWP U6922 ( .A1(n3579), .A2(\vrf/regTable[1][252] ), .B1(n7114), .B2(
        \vrf/regTable[3][252] ), .ZN(n8112) );
  AOI22D1BWP U6923 ( .A1(n8278), .A2(\vrf/regTable[0][252] ), .B1(n7110), .B2(
        \vrf/regTable[2][252] ), .ZN(n8111) );
  AOI211XD0BWP U6924 ( .A1(n5228), .A2(vectorData1[220]), .B(n5099), .C(n5098), 
        .ZN(n5100) );
  ND4D1BWP U6925 ( .A1(n5097), .A2(n5096), .A3(n5095), .A4(n5094), .ZN(n5098)
         );
  AOI22D1BWP U6926 ( .A1(n5231), .A2(vectorData1[124]), .B1(n5186), .B2(
        vectorData1[76]), .ZN(n5094) );
  ND4D1BWP U6927 ( .A1(n7407), .A2(n7408), .A3(n7409), .A4(n7410), .ZN(
        vectorData1[76]) );
  AOI22D1BWP U6928 ( .A1(n3576), .A2(\vrf/regTable[5][76] ), .B1(n3567), .B2(
        \vrf/regTable[7][76] ), .ZN(n7410) );
  AOI22D1BWP U6929 ( .A1(n3574), .A2(\vrf/regTable[4][76] ), .B1(n3570), .B2(
        \vrf/regTable[6][76] ), .ZN(n7409) );
  AOI22D1BWP U6930 ( .A1(n3579), .A2(\vrf/regTable[1][76] ), .B1(n3575), .B2(
        \vrf/regTable[3][76] ), .ZN(n7408) );
  AOI22D1BWP U6931 ( .A1(n3581), .A2(\vrf/regTable[0][76] ), .B1(n3572), .B2(
        \vrf/regTable[2][76] ), .ZN(n7407) );
  ND4D1BWP U6932 ( .A1(n7599), .A2(n7600), .A3(n7601), .A4(n7602), .ZN(
        vectorData1[124]) );
  AOI22D1BWP U6933 ( .A1(n7117), .A2(\vrf/regTable[5][124] ), .B1(n3567), .B2(
        \vrf/regTable[7][124] ), .ZN(n7602) );
  AOI22D1BWP U6934 ( .A1(n7115), .A2(\vrf/regTable[4][124] ), .B1(n3570), .B2(
        \vrf/regTable[6][124] ), .ZN(n7601) );
  AOI22D1BWP U6935 ( .A1(n7112), .A2(\vrf/regTable[1][124] ), .B1(n3599), .B2(
        \vrf/regTable[3][124] ), .ZN(n7600) );
  AOI22D1BWP U6936 ( .A1(n7108), .A2(\vrf/regTable[0][124] ), .B1(n3572), .B2(
        \vrf/regTable[2][124] ), .ZN(n7599) );
  AOI22D1BWP U6937 ( .A1(n5187), .A2(vectorData1[236]), .B1(n5188), .B2(
        vectorData1[60]), .ZN(n5095) );
  ND4D1BWP U6938 ( .A1(n7343), .A2(n7344), .A3(n7345), .A4(n7346), .ZN(
        vectorData1[60]) );
  AOI22D1BWP U6939 ( .A1(n3576), .A2(\vrf/regTable[5][60] ), .B1(n3567), .B2(
        \vrf/regTable[7][60] ), .ZN(n7346) );
  AOI22D1BWP U6940 ( .A1(n7115), .A2(\vrf/regTable[4][60] ), .B1(n3570), .B2(
        \vrf/regTable[6][60] ), .ZN(n7345) );
  AOI22D1BWP U6941 ( .A1(n3579), .A2(\vrf/regTable[1][60] ), .B1(n3575), .B2(
        \vrf/regTable[3][60] ), .ZN(n7344) );
  AOI22D1BWP U6942 ( .A1(n7108), .A2(\vrf/regTable[0][60] ), .B1(n3572), .B2(
        \vrf/regTable[2][60] ), .ZN(n7343) );
  ND4D1BWP U6943 ( .A1(n8047), .A2(n8048), .A3(n8049), .A4(n8050), .ZN(
        vectorData1[236]) );
  AOI22D1BWP U6944 ( .A1(n3576), .A2(\vrf/regTable[5][236] ), .B1(n3595), .B2(
        \vrf/regTable[7][236] ), .ZN(n8050) );
  AOI22D1BWP U6945 ( .A1(n8285), .A2(\vrf/regTable[4][236] ), .B1(n3596), .B2(
        \vrf/regTable[6][236] ), .ZN(n8049) );
  AOI22D1BWP U6946 ( .A1(n3579), .A2(\vrf/regTable[1][236] ), .B1(n3599), .B2(
        \vrf/regTable[3][236] ), .ZN(n8048) );
  AOI22D1BWP U6947 ( .A1(n8278), .A2(\vrf/regTable[0][236] ), .B1(n3594), .B2(
        \vrf/regTable[2][236] ), .ZN(n8047) );
  AOI22D1BWP U6948 ( .A1(n5233), .A2(vectorData1[188]), .B1(n5232), .B2(
        vectorData1[156]), .ZN(n5096) );
  ND4D1BWP U6949 ( .A1(n7727), .A2(n7728), .A3(n7729), .A4(n7730), .ZN(
        vectorData1[156]) );
  AOI22D1BWP U6950 ( .A1(n3576), .A2(\vrf/regTable[5][156] ), .B1(n3567), .B2(
        \vrf/regTable[7][156] ), .ZN(n7730) );
  AOI22D1BWP U6951 ( .A1(n7115), .A2(\vrf/regTable[4][156] ), .B1(n3570), .B2(
        \vrf/regTable[6][156] ), .ZN(n7729) );
  AOI22D1BWP U6952 ( .A1(n3579), .A2(\vrf/regTable[1][156] ), .B1(n3599), .B2(
        \vrf/regTable[3][156] ), .ZN(n7728) );
  AOI22D1BWP U6953 ( .A1(n7108), .A2(\vrf/regTable[0][156] ), .B1(n3572), .B2(
        \vrf/regTable[2][156] ), .ZN(n7727) );
  ND4D1BWP U6954 ( .A1(n7855), .A2(n7856), .A3(n7857), .A4(n7858), .ZN(
        vectorData1[188]) );
  AOI22D1BWP U6955 ( .A1(n3576), .A2(\vrf/regTable[5][188] ), .B1(n3567), .B2(
        \vrf/regTable[7][188] ), .ZN(n7858) );
  AOI22D1BWP U6956 ( .A1(n3574), .A2(\vrf/regTable[4][188] ), .B1(n3570), .B2(
        \vrf/regTable[6][188] ), .ZN(n7857) );
  AOI22D1BWP U6957 ( .A1(n3579), .A2(\vrf/regTable[1][188] ), .B1(n3575), .B2(
        \vrf/regTable[3][188] ), .ZN(n7856) );
  AOI22D1BWP U6958 ( .A1(n3581), .A2(\vrf/regTable[0][188] ), .B1(n3572), .B2(
        \vrf/regTable[2][188] ), .ZN(n7855) );
  AOI22D1BWP U6959 ( .A1(n5213), .A2(vectorData1[108]), .B1(n5185), .B2(
        vectorData1[92]), .ZN(n5097) );
  ND4D1BWP U6960 ( .A1(n7471), .A2(n7472), .A3(n7473), .A4(n7474), .ZN(
        vectorData1[92]) );
  AOI22D1BWP U6961 ( .A1(n7117), .A2(\vrf/regTable[5][92] ), .B1(n3567), .B2(
        \vrf/regTable[7][92] ), .ZN(n7474) );
  AOI22D1BWP U6962 ( .A1(n7115), .A2(\vrf/regTable[4][92] ), .B1(n3570), .B2(
        \vrf/regTable[6][92] ), .ZN(n7473) );
  AOI22D1BWP U6963 ( .A1(n7112), .A2(\vrf/regTable[1][92] ), .B1(n3575), .B2(
        \vrf/regTable[3][92] ), .ZN(n7472) );
  AOI22D1BWP U6964 ( .A1(n7108), .A2(\vrf/regTable[0][92] ), .B1(n3572), .B2(
        \vrf/regTable[2][92] ), .ZN(n7471) );
  ND4D1BWP U6965 ( .A1(n7535), .A2(n7536), .A3(n7537), .A4(n7538), .ZN(
        vectorData1[108]) );
  AOI22D1BWP U6966 ( .A1(n3576), .A2(\vrf/regTable[5][108] ), .B1(n3595), .B2(
        \vrf/regTable[7][108] ), .ZN(n7538) );
  AOI22D1BWP U6967 ( .A1(n3574), .A2(\vrf/regTable[4][108] ), .B1(n3596), .B2(
        \vrf/regTable[6][108] ), .ZN(n7537) );
  AOI22D1BWP U6968 ( .A1(n3579), .A2(\vrf/regTable[1][108] ), .B1(n3599), .B2(
        \vrf/regTable[3][108] ), .ZN(n7536) );
  AOI22D1BWP U6969 ( .A1(n3581), .A2(\vrf/regTable[0][108] ), .B1(n3594), .B2(
        \vrf/regTable[2][108] ), .ZN(n7535) );
  AO22D1BWP U6970 ( .A1(n5184), .A2(vectorData1[28]), .B1(n5227), .B2(
        vectorData1[204]), .Z(n5099) );
  ND4D1BWP U6971 ( .A1(n7919), .A2(n7920), .A3(n7921), .A4(n7922), .ZN(
        vectorData1[204]) );
  AOI22D1BWP U6972 ( .A1(n3576), .A2(\vrf/regTable[5][204] ), .B1(n7118), .B2(
        \vrf/regTable[7][204] ), .ZN(n7922) );
  AOI22D1BWP U6973 ( .A1(n3574), .A2(\vrf/regTable[4][204] ), .B1(n7116), .B2(
        \vrf/regTable[6][204] ), .ZN(n7921) );
  AOI22D1BWP U6974 ( .A1(n3579), .A2(\vrf/regTable[1][204] ), .B1(n7114), .B2(
        \vrf/regTable[3][204] ), .ZN(n7920) );
  AOI22D1BWP U6975 ( .A1(n3581), .A2(\vrf/regTable[0][204] ), .B1(n7110), .B2(
        \vrf/regTable[2][204] ), .ZN(n7919) );
  ND4D1BWP U6976 ( .A1(n7215), .A2(n7216), .A3(n7217), .A4(n7218), .ZN(
        vectorData1[28]) );
  AOI22D1BWP U6977 ( .A1(n3576), .A2(\vrf/regTable[5][28] ), .B1(n3595), .B2(
        \vrf/regTable[7][28] ), .ZN(n7218) );
  AOI22D1BWP U6978 ( .A1(n3574), .A2(\vrf/regTable[4][28] ), .B1(n3596), .B2(
        \vrf/regTable[6][28] ), .ZN(n7217) );
  AOI22D1BWP U6979 ( .A1(n3579), .A2(\vrf/regTable[1][28] ), .B1(n3599), .B2(
        \vrf/regTable[3][28] ), .ZN(n7216) );
  AOI22D1BWP U6980 ( .A1(n3581), .A2(\vrf/regTable[0][28] ), .B1(n3594), .B2(
        \vrf/regTable[2][28] ), .ZN(n7215) );
  ND4D1BWP U6981 ( .A1(n7983), .A2(n7984), .A3(n7985), .A4(n7986), .ZN(
        vectorData1[220]) );
  AOI22D1BWP U6982 ( .A1(n3576), .A2(\vrf/regTable[5][220] ), .B1(n7118), .B2(
        \vrf/regTable[7][220] ), .ZN(n7986) );
  AOI22D1BWP U6983 ( .A1(n7115), .A2(\vrf/regTable[4][220] ), .B1(n7116), .B2(
        \vrf/regTable[6][220] ), .ZN(n7985) );
  AOI22D1BWP U6984 ( .A1(n3579), .A2(\vrf/regTable[1][220] ), .B1(n7114), .B2(
        \vrf/regTable[3][220] ), .ZN(n7984) );
  AOI22D1BWP U6985 ( .A1(n7108), .A2(\vrf/regTable[0][220] ), .B1(n7110), .B2(
        \vrf/regTable[2][220] ), .ZN(n7983) );
  AOI22D1BWP U6986 ( .A1(n5226), .A2(vectorData1[140]), .B1(n3601), .B2(
        vectorData1[44]), .ZN(n5101) );
  ND4D1BWP U6987 ( .A1(n7279), .A2(n7280), .A3(n7281), .A4(n7282), .ZN(
        vectorData1[44]) );
  AOI22D1BWP U6988 ( .A1(n3576), .A2(\vrf/regTable[5][44] ), .B1(n3595), .B2(
        \vrf/regTable[7][44] ), .ZN(n7282) );
  AOI22D1BWP U6989 ( .A1(n8285), .A2(\vrf/regTable[4][44] ), .B1(n3596), .B2(
        \vrf/regTable[6][44] ), .ZN(n7281) );
  AOI22D1BWP U6990 ( .A1(n3579), .A2(\vrf/regTable[1][44] ), .B1(n3599), .B2(
        \vrf/regTable[3][44] ), .ZN(n7280) );
  AOI22D1BWP U6991 ( .A1(n8278), .A2(\vrf/regTable[0][44] ), .B1(n3594), .B2(
        \vrf/regTable[2][44] ), .ZN(n7279) );
  ND4D1BWP U6992 ( .A1(n7663), .A2(n7664), .A3(n7665), .A4(n7666), .ZN(
        vectorData1[140]) );
  AOI22D1BWP U6993 ( .A1(n3576), .A2(\vrf/regTable[5][140] ), .B1(n3567), .B2(
        \vrf/regTable[7][140] ), .ZN(n7666) );
  AOI22D1BWP U6994 ( .A1(n3574), .A2(\vrf/regTable[4][140] ), .B1(n3570), .B2(
        \vrf/regTable[6][140] ), .ZN(n7665) );
  AOI22D1BWP U6995 ( .A1(n3579), .A2(\vrf/regTable[1][140] ), .B1(n3599), .B2(
        \vrf/regTable[3][140] ), .ZN(n7664) );
  AOI22D1BWP U6996 ( .A1(n3581), .A2(\vrf/regTable[0][140] ), .B1(n3572), .B2(
        \vrf/regTable[2][140] ), .ZN(n7663) );
  ND4D1BWP U6997 ( .A1(n8325), .A2(n8326), .A3(n8327), .A4(n8328), .ZN(
        scalarData1[12]) );
  AOI22D1BWP U6998 ( .A1(n8287), .A2(\srf/regTable[5][12] ), .B1(n8288), .B2(
        \srf/regTable[7][12] ), .ZN(n8328) );
  AOI22D1BWP U6999 ( .A1(n8285), .A2(\srf/regTable[4][12] ), .B1(n8286), .B2(
        \srf/regTable[6][12] ), .ZN(n8327) );
  AOI22D1BWP U7000 ( .A1(n8282), .A2(\srf/regTable[1][12] ), .B1(n8284), .B2(
        \srf/regTable[3][12] ), .ZN(n8326) );
  AOI22D1BWP U7001 ( .A1(n8278), .A2(\srf/regTable[0][12] ), .B1(n8280), .B2(
        \srf/regTable[2][12] ), .ZN(n8325) );
  OAI211D1BWP U7002 ( .A1(n5443), .A2(n4405), .B(n5319), .C(n4535), .ZN(N4355)
         );
  AOI22D1BWP U7003 ( .A1(result[9]), .A2(n5331), .B1(n3668), .B2(
        vectorToLoad[137]), .ZN(n5319) );
  OAI211D1BWP U7004 ( .A1(n5446), .A2(n4405), .B(n5321), .C(n4535), .ZN(N4356)
         );
  AOI22D1BWP U7005 ( .A1(result[10]), .A2(n5331), .B1(n3668), .B2(
        vectorToLoad[138]), .ZN(n5321) );
  AO222D1BWP U7006 ( .A1(n3668), .A2(vectorToLoad[53]), .B1(n5394), .B2(n3649), 
        .C1(n4549), .C2(n5543), .Z(N4270) );
  ND4D1BWP U7007 ( .A1(n8043), .A2(n8044), .A3(n8045), .A4(n8046), .ZN(
        vectorData1[235]) );
  AOI22D1BWP U7008 ( .A1(n3576), .A2(\vrf/regTable[5][235] ), .B1(n3595), .B2(
        \vrf/regTable[7][235] ), .ZN(n8046) );
  AOI22D1BWP U7009 ( .A1(n7115), .A2(\vrf/regTable[4][235] ), .B1(n3596), .B2(
        \vrf/regTable[6][235] ), .ZN(n8045) );
  AOI22D1BWP U7010 ( .A1(n3579), .A2(\vrf/regTable[1][235] ), .B1(n3599), .B2(
        \vrf/regTable[3][235] ), .ZN(n8044) );
  AOI22D1BWP U7011 ( .A1(n7108), .A2(\vrf/regTable[0][235] ), .B1(n3594), .B2(
        \vrf/regTable[2][235] ), .ZN(n8043) );
  ND4D1BWP U7012 ( .A1(n8107), .A2(n8108), .A3(n8109), .A4(n8110), .ZN(
        vectorData1[251]) );
  AOI22D1BWP U7013 ( .A1(n3576), .A2(\vrf/regTable[5][251] ), .B1(n7118), .B2(
        \vrf/regTable[7][251] ), .ZN(n8110) );
  AOI22D1BWP U7014 ( .A1(n3574), .A2(\vrf/regTable[4][251] ), .B1(n7116), .B2(
        \vrf/regTable[6][251] ), .ZN(n8109) );
  AOI22D1BWP U7015 ( .A1(n3579), .A2(\vrf/regTable[1][251] ), .B1(n7114), .B2(
        \vrf/regTable[3][251] ), .ZN(n8108) );
  AOI22D1BWP U7016 ( .A1(n3581), .A2(\vrf/regTable[0][251] ), .B1(n7110), .B2(
        \vrf/regTable[2][251] ), .ZN(n8107) );
  ND4D1BWP U7017 ( .A1(n5092), .A2(n5091), .A3(n5090), .A4(n5089), .ZN(n5093)
         );
  AOI22D1BWP U7018 ( .A1(n5185), .A2(vectorData1[91]), .B1(n5188), .B2(
        vectorData1[59]), .ZN(n5089) );
  ND4D1BWP U7019 ( .A1(n7339), .A2(n7340), .A3(n7341), .A4(n7342), .ZN(
        vectorData1[59]) );
  AOI22D1BWP U7020 ( .A1(n3576), .A2(\vrf/regTable[5][59] ), .B1(n3567), .B2(
        \vrf/regTable[7][59] ), .ZN(n7342) );
  AOI22D1BWP U7021 ( .A1(n3574), .A2(\vrf/regTable[4][59] ), .B1(n3570), .B2(
        \vrf/regTable[6][59] ), .ZN(n7341) );
  AOI22D1BWP U7022 ( .A1(n3579), .A2(\vrf/regTable[1][59] ), .B1(n3575), .B2(
        \vrf/regTable[3][59] ), .ZN(n7340) );
  AOI22D1BWP U7023 ( .A1(n3581), .A2(\vrf/regTable[0][59] ), .B1(n3572), .B2(
        \vrf/regTable[2][59] ), .ZN(n7339) );
  ND4D1BWP U7024 ( .A1(n7467), .A2(n7468), .A3(n7469), .A4(n7470), .ZN(
        vectorData1[91]) );
  AOI22D1BWP U7025 ( .A1(n3576), .A2(\vrf/regTable[5][91] ), .B1(n3567), .B2(
        \vrf/regTable[7][91] ), .ZN(n7470) );
  AOI22D1BWP U7026 ( .A1(n8285), .A2(\vrf/regTable[4][91] ), .B1(n3570), .B2(
        \vrf/regTable[6][91] ), .ZN(n7469) );
  AOI22D1BWP U7027 ( .A1(n3579), .A2(\vrf/regTable[1][91] ), .B1(n3575), .B2(
        \vrf/regTable[3][91] ), .ZN(n7468) );
  AOI22D1BWP U7028 ( .A1(n8278), .A2(\vrf/regTable[0][91] ), .B1(n3572), .B2(
        \vrf/regTable[2][91] ), .ZN(n7467) );
  AOI22D1BWP U7029 ( .A1(n5184), .A2(vectorData1[27]), .B1(n5227), .B2(
        vectorData1[203]), .ZN(n5090) );
  ND4D1BWP U7030 ( .A1(n7915), .A2(n7916), .A3(n7917), .A4(n7918), .ZN(
        vectorData1[203]) );
  AOI22D1BWP U7031 ( .A1(n3576), .A2(\vrf/regTable[5][203] ), .B1(n3595), .B2(
        \vrf/regTable[7][203] ), .ZN(n7918) );
  AOI22D1BWP U7032 ( .A1(n3574), .A2(\vrf/regTable[4][203] ), .B1(n3596), .B2(
        \vrf/regTable[6][203] ), .ZN(n7917) );
  AOI22D1BWP U7033 ( .A1(n3579), .A2(\vrf/regTable[1][203] ), .B1(n3599), .B2(
        \vrf/regTable[3][203] ), .ZN(n7916) );
  AOI22D1BWP U7034 ( .A1(n3581), .A2(\vrf/regTable[0][203] ), .B1(n3594), .B2(
        \vrf/regTable[2][203] ), .ZN(n7915) );
  ND4D1BWP U7035 ( .A1(n7211), .A2(n7212), .A3(n7213), .A4(n7214), .ZN(
        vectorData1[27]) );
  AOI22D1BWP U7036 ( .A1(n3576), .A2(\vrf/regTable[5][27] ), .B1(n3595), .B2(
        \vrf/regTable[7][27] ), .ZN(n7214) );
  AOI22D1BWP U7037 ( .A1(n7115), .A2(\vrf/regTable[4][27] ), .B1(n3596), .B2(
        \vrf/regTable[6][27] ), .ZN(n7213) );
  AOI22D1BWP U7038 ( .A1(n3579), .A2(\vrf/regTable[1][27] ), .B1(n3599), .B2(
        \vrf/regTable[3][27] ), .ZN(n7212) );
  AOI22D1BWP U7039 ( .A1(n7108), .A2(\vrf/regTable[0][27] ), .B1(n3594), .B2(
        \vrf/regTable[2][27] ), .ZN(n7211) );
  AOI22D1BWP U7040 ( .A1(n5228), .A2(vectorData1[219]), .B1(n5230), .B2(
        vectorData1[171]), .ZN(n5091) );
  ND4D1BWP U7041 ( .A1(n7787), .A2(n7788), .A3(n7789), .A4(n7790), .ZN(
        vectorData1[171]) );
  AOI22D1BWP U7042 ( .A1(n3576), .A2(\vrf/regTable[5][171] ), .B1(n3567), .B2(
        \vrf/regTable[7][171] ), .ZN(n7790) );
  AOI22D1BWP U7043 ( .A1(n8285), .A2(\vrf/regTable[4][171] ), .B1(n3570), .B2(
        \vrf/regTable[6][171] ), .ZN(n7789) );
  AOI22D1BWP U7044 ( .A1(n3579), .A2(\vrf/regTable[1][171] ), .B1(n3575), .B2(
        \vrf/regTable[3][171] ), .ZN(n7788) );
  AOI22D1BWP U7045 ( .A1(n8278), .A2(\vrf/regTable[0][171] ), .B1(n3572), .B2(
        \vrf/regTable[2][171] ), .ZN(n7787) );
  ND4D1BWP U7046 ( .A1(n7979), .A2(n7980), .A3(n7981), .A4(n7982), .ZN(
        vectorData1[219]) );
  AOI22D1BWP U7047 ( .A1(n3576), .A2(\vrf/regTable[5][219] ), .B1(n3567), .B2(
        \vrf/regTable[7][219] ), .ZN(n7982) );
  AOI22D1BWP U7048 ( .A1(n3574), .A2(\vrf/regTable[4][219] ), .B1(n3570), .B2(
        \vrf/regTable[6][219] ), .ZN(n7981) );
  AOI22D1BWP U7049 ( .A1(n3579), .A2(\vrf/regTable[1][219] ), .B1(n3575), .B2(
        \vrf/regTable[3][219] ), .ZN(n7980) );
  AOI22D1BWP U7050 ( .A1(n3581), .A2(\vrf/regTable[0][219] ), .B1(n3572), .B2(
        \vrf/regTable[2][219] ), .ZN(n7979) );
  AOI22D1BWP U7051 ( .A1(n5233), .A2(vectorData1[187]), .B1(n3601), .B2(
        vectorData1[43]), .ZN(n5092) );
  ND4D1BWP U7052 ( .A1(n7275), .A2(n7276), .A3(n7277), .A4(n7278), .ZN(
        vectorData1[43]) );
  AOI22D1BWP U7053 ( .A1(n3576), .A2(\vrf/regTable[5][43] ), .B1(n3595), .B2(
        \vrf/regTable[7][43] ), .ZN(n7278) );
  AOI22D1BWP U7054 ( .A1(n3574), .A2(\vrf/regTable[4][43] ), .B1(n3596), .B2(
        \vrf/regTable[6][43] ), .ZN(n7277) );
  AOI22D1BWP U7055 ( .A1(n3579), .A2(\vrf/regTable[1][43] ), .B1(n3599), .B2(
        \vrf/regTable[3][43] ), .ZN(n7276) );
  AOI22D1BWP U7056 ( .A1(n3581), .A2(\vrf/regTable[0][43] ), .B1(n3594), .B2(
        \vrf/regTable[2][43] ), .ZN(n7275) );
  ND4D1BWP U7057 ( .A1(n7851), .A2(n7852), .A3(n7853), .A4(n7854), .ZN(
        vectorData1[187]) );
  AOI22D1BWP U7058 ( .A1(n3576), .A2(\vrf/regTable[5][187] ), .B1(n3567), .B2(
        \vrf/regTable[7][187] ), .ZN(n7854) );
  AOI22D1BWP U7059 ( .A1(n3574), .A2(\vrf/regTable[4][187] ), .B1(n3570), .B2(
        \vrf/regTable[6][187] ), .ZN(n7853) );
  AOI22D1BWP U7060 ( .A1(n3579), .A2(\vrf/regTable[1][187] ), .B1(n3575), .B2(
        \vrf/regTable[3][187] ), .ZN(n7852) );
  AOI22D1BWP U7061 ( .A1(n3581), .A2(\vrf/regTable[0][187] ), .B1(n3572), .B2(
        \vrf/regTable[2][187] ), .ZN(n7851) );
  ND4D1BWP U7062 ( .A1(n7723), .A2(n7724), .A3(n7725), .A4(n7726), .ZN(
        vectorData1[155]) );
  AOI22D1BWP U7063 ( .A1(n3576), .A2(\vrf/regTable[5][155] ), .B1(n3595), .B2(
        \vrf/regTable[7][155] ), .ZN(n7726) );
  AOI22D1BWP U7064 ( .A1(n3574), .A2(\vrf/regTable[4][155] ), .B1(n3596), .B2(
        \vrf/regTable[6][155] ), .ZN(n7725) );
  AOI22D1BWP U7065 ( .A1(n3579), .A2(\vrf/regTable[1][155] ), .B1(n3575), .B2(
        \vrf/regTable[3][155] ), .ZN(n7724) );
  AOI22D1BWP U7066 ( .A1(n3581), .A2(\vrf/regTable[0][155] ), .B1(n3594), .B2(
        \vrf/regTable[2][155] ), .ZN(n7723) );
  ND4D1BWP U7067 ( .A1(n7531), .A2(n7532), .A3(n7533), .A4(n7534), .ZN(
        vectorData1[107]) );
  AOI22D1BWP U7068 ( .A1(n3576), .A2(\vrf/regTable[5][107] ), .B1(n3595), .B2(
        \vrf/regTable[7][107] ), .ZN(n7534) );
  AOI22D1BWP U7069 ( .A1(n3574), .A2(\vrf/regTable[4][107] ), .B1(n3596), .B2(
        \vrf/regTable[6][107] ), .ZN(n7533) );
  AOI22D1BWP U7070 ( .A1(n3579), .A2(\vrf/regTable[1][107] ), .B1(n3575), .B2(
        \vrf/regTable[3][107] ), .ZN(n7532) );
  AOI22D1BWP U7071 ( .A1(n3581), .A2(\vrf/regTable[0][107] ), .B1(n3594), .B2(
        \vrf/regTable[2][107] ), .ZN(n7531) );
  ND4D1BWP U7072 ( .A1(n7659), .A2(n7660), .A3(n7661), .A4(n7662), .ZN(
        vectorData1[139]) );
  AOI22D1BWP U7073 ( .A1(n3576), .A2(\vrf/regTable[5][139] ), .B1(n3567), .B2(
        \vrf/regTable[7][139] ), .ZN(n7662) );
  AOI22D1BWP U7074 ( .A1(n3574), .A2(\vrf/regTable[4][139] ), .B1(n3570), .B2(
        \vrf/regTable[6][139] ), .ZN(n7661) );
  AOI22D1BWP U7075 ( .A1(n3579), .A2(\vrf/regTable[1][139] ), .B1(n3599), .B2(
        \vrf/regTable[3][139] ), .ZN(n7660) );
  AOI22D1BWP U7076 ( .A1(n3581), .A2(\vrf/regTable[0][139] ), .B1(n3572), .B2(
        \vrf/regTable[2][139] ), .ZN(n7659) );
  AOI22D1BWP U7077 ( .A1(n3576), .A2(\vrf/regTable[5][75] ), .B1(n3595), .B2(
        \vrf/regTable[7][75] ), .ZN(n7406) );
  AOI22D1BWP U7078 ( .A1(n3574), .A2(\vrf/regTable[4][75] ), .B1(n3596), .B2(
        \vrf/regTable[6][75] ), .ZN(n7405) );
  AOI22D1BWP U7079 ( .A1(n3579), .A2(\vrf/regTable[1][75] ), .B1(n3599), .B2(
        \vrf/regTable[3][75] ), .ZN(n7404) );
  AOI22D1BWP U7080 ( .A1(n3581), .A2(\vrf/regTable[0][75] ), .B1(n3594), .B2(
        \vrf/regTable[2][75] ), .ZN(n7403) );
  AOI22D1BWP U7081 ( .A1(n3576), .A2(\vrf/regTable[5][123] ), .B1(n3567), .B2(
        \vrf/regTable[7][123] ), .ZN(n7598) );
  AOI22D1BWP U7082 ( .A1(n3574), .A2(\vrf/regTable[4][123] ), .B1(n3570), .B2(
        \vrf/regTable[6][123] ), .ZN(n7597) );
  AOI22D1BWP U7083 ( .A1(n3579), .A2(\vrf/regTable[1][123] ), .B1(n3599), .B2(
        \vrf/regTable[3][123] ), .ZN(n7596) );
  AOI22D1BWP U7084 ( .A1(n3581), .A2(\vrf/regTable[0][123] ), .B1(n3572), .B2(
        \vrf/regTable[2][123] ), .ZN(n7595) );
  OAI211D1BWP U7085 ( .A1(n5449), .A2(n4405), .B(n5323), .C(n4535), .ZN(N4357)
         );
  AOI22D1BWP U7086 ( .A1(result[11]), .A2(n5331), .B1(n3668), .B2(
        vectorToLoad[139]), .ZN(n5323) );
  AO222D1BWP U7087 ( .A1(n3639), .A2(n4548), .B1(n5525), .B2(n4628), .C1(n4631), .C2(vectorToLoad[101]), .Z(N4318) );
  OAI211D1BWP U7088 ( .A1(n5452), .A2(n4405), .B(n5325), .C(n4535), .ZN(N4358)
         );
  AOI22D1BWP U7089 ( .A1(result[12]), .A2(n5331), .B1(n3668), .B2(
        vectorToLoad[140]), .ZN(n5325) );
  ND4D1BWP U7090 ( .A1(n7719), .A2(n7720), .A3(n7721), .A4(n7722), .ZN(
        vectorData1[154]) );
  AOI22D1BWP U7091 ( .A1(n3576), .A2(\vrf/regTable[5][154] ), .B1(n3567), .B2(
        \vrf/regTable[7][154] ), .ZN(n7722) );
  AOI22D1BWP U7092 ( .A1(n3574), .A2(\vrf/regTable[4][154] ), .B1(n3570), .B2(
        \vrf/regTable[6][154] ), .ZN(n7721) );
  AOI22D1BWP U7093 ( .A1(n3579), .A2(\vrf/regTable[1][154] ), .B1(n3599), .B2(
        \vrf/regTable[3][154] ), .ZN(n7720) );
  AOI22D1BWP U7094 ( .A1(n3581), .A2(\vrf/regTable[0][154] ), .B1(n3572), .B2(
        \vrf/regTable[2][154] ), .ZN(n7719) );
  ND4D1BWP U7095 ( .A1(n7463), .A2(n7464), .A3(n7465), .A4(n7466), .ZN(
        vectorData1[90]) );
  AOI22D1BWP U7096 ( .A1(n7117), .A2(\vrf/regTable[5][90] ), .B1(n3567), .B2(
        \vrf/regTable[7][90] ), .ZN(n7466) );
  AOI22D1BWP U7097 ( .A1(n7115), .A2(\vrf/regTable[4][90] ), .B1(n3570), .B2(
        \vrf/regTable[6][90] ), .ZN(n7465) );
  AOI22D1BWP U7098 ( .A1(n7112), .A2(\vrf/regTable[1][90] ), .B1(n3575), .B2(
        \vrf/regTable[3][90] ), .ZN(n7464) );
  AOI22D1BWP U7099 ( .A1(n7108), .A2(\vrf/regTable[0][90] ), .B1(n3572), .B2(
        \vrf/regTable[2][90] ), .ZN(n7463) );
  ND4D1BWP U7100 ( .A1(n5087), .A2(n5086), .A3(n5085), .A4(n5084), .ZN(n5088)
         );
  AOI22D1BWP U7101 ( .A1(n5226), .A2(vectorData1[138]), .B1(n5229), .B2(
        vectorData1[250]), .ZN(n5084) );
  ND4D1BWP U7102 ( .A1(n8103), .A2(n8104), .A3(n8105), .A4(n8106), .ZN(
        vectorData1[250]) );
  AOI22D1BWP U7103 ( .A1(n3576), .A2(\vrf/regTable[5][250] ), .B1(n3595), .B2(
        \vrf/regTable[7][250] ), .ZN(n8106) );
  AOI22D1BWP U7104 ( .A1(n3574), .A2(\vrf/regTable[4][250] ), .B1(n3596), .B2(
        \vrf/regTable[6][250] ), .ZN(n8105) );
  AOI22D1BWP U7105 ( .A1(n3579), .A2(\vrf/regTable[1][250] ), .B1(n3599), .B2(
        \vrf/regTable[3][250] ), .ZN(n8104) );
  AOI22D1BWP U7106 ( .A1(n3581), .A2(\vrf/regTable[0][250] ), .B1(n3594), .B2(
        \vrf/regTable[2][250] ), .ZN(n8103) );
  ND4D1BWP U7107 ( .A1(n7655), .A2(n7656), .A3(n7657), .A4(n7658), .ZN(
        vectorData1[138]) );
  AOI22D1BWP U7108 ( .A1(n3576), .A2(\vrf/regTable[5][138] ), .B1(n3567), .B2(
        \vrf/regTable[7][138] ), .ZN(n7658) );
  AOI22D1BWP U7109 ( .A1(n3574), .A2(\vrf/regTable[4][138] ), .B1(n3570), .B2(
        \vrf/regTable[6][138] ), .ZN(n7657) );
  AOI22D1BWP U7110 ( .A1(n3579), .A2(\vrf/regTable[1][138] ), .B1(n3599), .B2(
        \vrf/regTable[3][138] ), .ZN(n7656) );
  AOI22D1BWP U7111 ( .A1(n3581), .A2(\vrf/regTable[0][138] ), .B1(n3572), .B2(
        \vrf/regTable[2][138] ), .ZN(n7655) );
  AOI22D1BWP U7112 ( .A1(n5228), .A2(vectorData1[218]), .B1(n5187), .B2(
        vectorData1[234]), .ZN(n5085) );
  ND4D1BWP U7113 ( .A1(n8039), .A2(n8040), .A3(n8041), .A4(n8042), .ZN(
        vectorData1[234]) );
  AOI22D1BWP U7114 ( .A1(n3576), .A2(\vrf/regTable[5][234] ), .B1(n7118), .B2(
        \vrf/regTable[7][234] ), .ZN(n8042) );
  AOI22D1BWP U7115 ( .A1(n7115), .A2(\vrf/regTable[4][234] ), .B1(n7116), .B2(
        \vrf/regTable[6][234] ), .ZN(n8041) );
  AOI22D1BWP U7116 ( .A1(n3579), .A2(\vrf/regTable[1][234] ), .B1(n7114), .B2(
        \vrf/regTable[3][234] ), .ZN(n8040) );
  AOI22D1BWP U7117 ( .A1(n7108), .A2(\vrf/regTable[0][234] ), .B1(n7110), .B2(
        \vrf/regTable[2][234] ), .ZN(n8039) );
  ND4D1BWP U7118 ( .A1(n7975), .A2(n7976), .A3(n7977), .A4(n7978), .ZN(
        vectorData1[218]) );
  AOI22D1BWP U7119 ( .A1(n3576), .A2(\vrf/regTable[5][218] ), .B1(n3595), .B2(
        \vrf/regTable[7][218] ), .ZN(n7978) );
  AOI22D1BWP U7120 ( .A1(n3574), .A2(\vrf/regTable[4][218] ), .B1(n3596), .B2(
        \vrf/regTable[6][218] ), .ZN(n7977) );
  AOI22D1BWP U7121 ( .A1(n3579), .A2(\vrf/regTable[1][218] ), .B1(n3599), .B2(
        \vrf/regTable[3][218] ), .ZN(n7976) );
  AOI22D1BWP U7122 ( .A1(n3581), .A2(\vrf/regTable[0][218] ), .B1(n3594), .B2(
        \vrf/regTable[2][218] ), .ZN(n7975) );
  AOI22D1BWP U7123 ( .A1(n5231), .A2(vectorData1[122]), .B1(n5227), .B2(
        vectorData1[202]), .ZN(n5086) );
  ND4D1BWP U7124 ( .A1(n7911), .A2(n7912), .A3(n7913), .A4(n7914), .ZN(
        vectorData1[202]) );
  AOI22D1BWP U7125 ( .A1(n3576), .A2(\vrf/regTable[5][202] ), .B1(n3595), .B2(
        \vrf/regTable[7][202] ), .ZN(n7914) );
  AOI22D1BWP U7126 ( .A1(n3574), .A2(\vrf/regTable[4][202] ), .B1(n3596), .B2(
        \vrf/regTable[6][202] ), .ZN(n7913) );
  AOI22D1BWP U7127 ( .A1(n3579), .A2(\vrf/regTable[1][202] ), .B1(n3599), .B2(
        \vrf/regTable[3][202] ), .ZN(n7912) );
  AOI22D1BWP U7128 ( .A1(n3581), .A2(\vrf/regTable[0][202] ), .B1(n3594), .B2(
        \vrf/regTable[2][202] ), .ZN(n7911) );
  ND4D1BWP U7129 ( .A1(n7591), .A2(n7592), .A3(n7593), .A4(n7594), .ZN(
        vectorData1[122]) );
  AOI22D1BWP U7130 ( .A1(n3576), .A2(\vrf/regTable[5][122] ), .B1(n3595), .B2(
        \vrf/regTable[7][122] ), .ZN(n7594) );
  AOI22D1BWP U7131 ( .A1(n3574), .A2(\vrf/regTable[4][122] ), .B1(n3596), .B2(
        \vrf/regTable[6][122] ), .ZN(n7593) );
  AOI22D1BWP U7132 ( .A1(n3579), .A2(\vrf/regTable[1][122] ), .B1(n3575), .B2(
        \vrf/regTable[3][122] ), .ZN(n7592) );
  AOI22D1BWP U7133 ( .A1(n3581), .A2(\vrf/regTable[0][122] ), .B1(n3594), .B2(
        \vrf/regTable[2][122] ), .ZN(n7591) );
  AOI22D1BWP U7134 ( .A1(n5184), .A2(vectorData1[26]), .B1(n5186), .B2(
        vectorData1[74]), .ZN(n5087) );
  ND4D1BWP U7135 ( .A1(n7399), .A2(n7400), .A3(n7401), .A4(n7402), .ZN(
        vectorData1[74]) );
  AOI22D1BWP U7136 ( .A1(n3576), .A2(\vrf/regTable[5][74] ), .B1(n3567), .B2(
        \vrf/regTable[7][74] ), .ZN(n7402) );
  AOI22D1BWP U7137 ( .A1(n8285), .A2(\vrf/regTable[4][74] ), .B1(n3570), .B2(
        \vrf/regTable[6][74] ), .ZN(n7401) );
  AOI22D1BWP U7138 ( .A1(n3579), .A2(\vrf/regTable[1][74] ), .B1(n3575), .B2(
        \vrf/regTable[3][74] ), .ZN(n7400) );
  AOI22D1BWP U7139 ( .A1(n8278), .A2(\vrf/regTable[0][74] ), .B1(n3572), .B2(
        \vrf/regTable[2][74] ), .ZN(n7399) );
  ND4D1BWP U7140 ( .A1(n7207), .A2(n7208), .A3(n7209), .A4(n7210), .ZN(
        vectorData1[26]) );
  AOI22D1BWP U7141 ( .A1(n3576), .A2(\vrf/regTable[5][26] ), .B1(n3567), .B2(
        \vrf/regTable[7][26] ), .ZN(n7210) );
  AOI22D1BWP U7142 ( .A1(n7115), .A2(\vrf/regTable[4][26] ), .B1(n3570), .B2(
        \vrf/regTable[6][26] ), .ZN(n7209) );
  AOI22D1BWP U7143 ( .A1(n3579), .A2(\vrf/regTable[1][26] ), .B1(n3575), .B2(
        \vrf/regTable[3][26] ), .ZN(n7208) );
  AOI22D1BWP U7144 ( .A1(n7108), .A2(\vrf/regTable[0][26] ), .B1(n3572), .B2(
        \vrf/regTable[2][26] ), .ZN(n7207) );
  ND4D1BWP U7145 ( .A1(n7783), .A2(n7784), .A3(n7785), .A4(n7786), .ZN(
        vectorData1[170]) );
  AOI22D1BWP U7146 ( .A1(n3576), .A2(\vrf/regTable[5][170] ), .B1(n3595), .B2(
        \vrf/regTable[7][170] ), .ZN(n7786) );
  AOI22D1BWP U7147 ( .A1(n7115), .A2(\vrf/regTable[4][170] ), .B1(n3596), .B2(
        \vrf/regTable[6][170] ), .ZN(n7785) );
  AOI22D1BWP U7148 ( .A1(n3579), .A2(\vrf/regTable[1][170] ), .B1(n3575), .B2(
        \vrf/regTable[3][170] ), .ZN(n7784) );
  AOI22D1BWP U7149 ( .A1(n7108), .A2(\vrf/regTable[0][170] ), .B1(n3594), .B2(
        \vrf/regTable[2][170] ), .ZN(n7783) );
  ND4D1BWP U7150 ( .A1(n7271), .A2(n7272), .A3(n7273), .A4(n7274), .ZN(
        vectorData1[42]) );
  AOI22D1BWP U7151 ( .A1(n3576), .A2(\vrf/regTable[5][42] ), .B1(n3595), .B2(
        \vrf/regTable[7][42] ), .ZN(n7274) );
  AOI22D1BWP U7152 ( .A1(n3574), .A2(\vrf/regTable[4][42] ), .B1(n3596), .B2(
        \vrf/regTable[6][42] ), .ZN(n7273) );
  AOI22D1BWP U7153 ( .A1(n3579), .A2(\vrf/regTable[1][42] ), .B1(n3599), .B2(
        \vrf/regTable[3][42] ), .ZN(n7272) );
  AOI22D1BWP U7154 ( .A1(n3581), .A2(\vrf/regTable[0][42] ), .B1(n3594), .B2(
        \vrf/regTable[2][42] ), .ZN(n7271) );
  ND4D1BWP U7155 ( .A1(n7847), .A2(n7848), .A3(n7849), .A4(n7850), .ZN(
        vectorData1[186]) );
  AOI22D1BWP U7156 ( .A1(n3576), .A2(\vrf/regTable[5][186] ), .B1(n3567), .B2(
        \vrf/regTable[7][186] ), .ZN(n7850) );
  AOI22D1BWP U7157 ( .A1(n3574), .A2(\vrf/regTable[4][186] ), .B1(n3570), .B2(
        \vrf/regTable[6][186] ), .ZN(n7849) );
  AOI22D1BWP U7158 ( .A1(n3579), .A2(\vrf/regTable[1][186] ), .B1(n3575), .B2(
        \vrf/regTable[3][186] ), .ZN(n7848) );
  AOI22D1BWP U7159 ( .A1(n3581), .A2(\vrf/regTable[0][186] ), .B1(n3572), .B2(
        \vrf/regTable[2][186] ), .ZN(n7847) );
  AOI22D1BWP U7160 ( .A1(n3576), .A2(\vrf/regTable[5][58] ), .B1(n3567), .B2(
        \vrf/regTable[7][58] ), .ZN(n7338) );
  AOI22D1BWP U7161 ( .A1(n3574), .A2(\vrf/regTable[4][58] ), .B1(n3570), .B2(
        \vrf/regTable[6][58] ), .ZN(n7337) );
  AOI22D1BWP U7162 ( .A1(n3579), .A2(\vrf/regTable[1][58] ), .B1(n3575), .B2(
        \vrf/regTable[3][58] ), .ZN(n7336) );
  AOI22D1BWP U7163 ( .A1(n3581), .A2(\vrf/regTable[0][58] ), .B1(n3572), .B2(
        \vrf/regTable[2][58] ), .ZN(n7335) );
  AOI22D1BWP U7164 ( .A1(n3576), .A2(\vrf/regTable[5][106] ), .B1(n3595), .B2(
        \vrf/regTable[7][106] ), .ZN(n7530) );
  AOI22D1BWP U7165 ( .A1(n3574), .A2(\vrf/regTable[4][106] ), .B1(n3596), .B2(
        \vrf/regTable[6][106] ), .ZN(n7529) );
  AOI22D1BWP U7166 ( .A1(n3579), .A2(\vrf/regTable[1][106] ), .B1(n3599), .B2(
        \vrf/regTable[3][106] ), .ZN(n7528) );
  AOI22D1BWP U7167 ( .A1(n3581), .A2(\vrf/regTable[0][106] ), .B1(n3594), .B2(
        \vrf/regTable[2][106] ), .ZN(n7527) );
  OAI211D1BWP U7168 ( .A1(n5455), .A2(n4405), .B(n5327), .C(n4535), .ZN(N4359)
         );
  AOI22D1BWP U7169 ( .A1(result[13]), .A2(n5331), .B1(n3668), .B2(
        vectorToLoad[141]), .ZN(n5327) );
  AO222D1BWP U7170 ( .A1(n3669), .A2(vectorToLoad[52]), .B1(n5341), .B2(n3649), 
        .C1(n4549), .C2(n5542), .Z(N4269) );
  OAI211D1BWP U7171 ( .A1(n5458), .A2(n4405), .B(n5329), .C(n4535), .ZN(N4360)
         );
  AOI22D1BWP U7172 ( .A1(result[14]), .A2(n5331), .B1(n3668), .B2(
        vectorToLoad[142]), .ZN(n5329) );
  ND4D1BWP U7173 ( .A1(n7907), .A2(n7908), .A3(n7909), .A4(n7910), .ZN(
        vectorData1[201]) );
  AOI22D1BWP U7174 ( .A1(n3576), .A2(\vrf/regTable[5][201] ), .B1(n3567), .B2(
        \vrf/regTable[7][201] ), .ZN(n7910) );
  AOI22D1BWP U7175 ( .A1(n3574), .A2(\vrf/regTable[4][201] ), .B1(n3570), .B2(
        \vrf/regTable[6][201] ), .ZN(n7909) );
  AOI22D1BWP U7176 ( .A1(n3579), .A2(\vrf/regTable[1][201] ), .B1(n3575), .B2(
        \vrf/regTable[3][201] ), .ZN(n7908) );
  AOI22D1BWP U7177 ( .A1(n3581), .A2(\vrf/regTable[0][201] ), .B1(n3572), .B2(
        \vrf/regTable[2][201] ), .ZN(n7907) );
  ND4D1BWP U7178 ( .A1(n8035), .A2(n8036), .A3(n8037), .A4(n8038), .ZN(
        vectorData1[233]) );
  AOI22D1BWP U7179 ( .A1(n3576), .A2(\vrf/regTable[5][233] ), .B1(n3595), .B2(
        \vrf/regTable[7][233] ), .ZN(n8038) );
  AOI22D1BWP U7180 ( .A1(n8285), .A2(\vrf/regTable[4][233] ), .B1(n3596), .B2(
        \vrf/regTable[6][233] ), .ZN(n8037) );
  AOI22D1BWP U7181 ( .A1(n3579), .A2(\vrf/regTable[1][233] ), .B1(n3599), .B2(
        \vrf/regTable[3][233] ), .ZN(n8036) );
  AOI22D1BWP U7182 ( .A1(n8278), .A2(\vrf/regTable[0][233] ), .B1(n3594), .B2(
        \vrf/regTable[2][233] ), .ZN(n8035) );
  AOI22D1BWP U7183 ( .A1(n5226), .A2(vectorData1[137]), .B1(n3601), .B2(
        vectorData1[41]), .ZN(n5080) );
  ND4D1BWP U7184 ( .A1(n7267), .A2(n7268), .A3(n7269), .A4(n7270), .ZN(
        vectorData1[41]) );
  AOI22D1BWP U7185 ( .A1(n3576), .A2(\vrf/regTable[5][41] ), .B1(n3595), .B2(
        \vrf/regTable[7][41] ), .ZN(n7270) );
  AOI22D1BWP U7186 ( .A1(n3574), .A2(\vrf/regTable[4][41] ), .B1(n3596), .B2(
        \vrf/regTable[6][41] ), .ZN(n7269) );
  AOI22D1BWP U7187 ( .A1(n3579), .A2(\vrf/regTable[1][41] ), .B1(n3599), .B2(
        \vrf/regTable[3][41] ), .ZN(n7268) );
  AOI22D1BWP U7188 ( .A1(n3581), .A2(\vrf/regTable[0][41] ), .B1(n3594), .B2(
        \vrf/regTable[2][41] ), .ZN(n7267) );
  ND4D1BWP U7189 ( .A1(n7651), .A2(n7652), .A3(n7653), .A4(n7654), .ZN(
        vectorData1[137]) );
  AOI22D1BWP U7190 ( .A1(n3576), .A2(\vrf/regTable[5][137] ), .B1(n3595), .B2(
        \vrf/regTable[7][137] ), .ZN(n7654) );
  AOI22D1BWP U7191 ( .A1(n7115), .A2(\vrf/regTable[4][137] ), .B1(n3596), .B2(
        \vrf/regTable[6][137] ), .ZN(n7653) );
  AOI22D1BWP U7192 ( .A1(n3579), .A2(\vrf/regTable[1][137] ), .B1(n3599), .B2(
        \vrf/regTable[3][137] ), .ZN(n7652) );
  AOI22D1BWP U7193 ( .A1(n7108), .A2(\vrf/regTable[0][137] ), .B1(n3594), .B2(
        \vrf/regTable[2][137] ), .ZN(n7651) );
  AOI22D1BWP U7194 ( .A1(n5228), .A2(vectorData1[217]), .B1(n5186), .B2(
        vectorData1[73]), .ZN(n5081) );
  ND4D1BWP U7195 ( .A1(n7395), .A2(n7396), .A3(n7397), .A4(n7398), .ZN(
        vectorData1[73]) );
  AOI22D1BWP U7196 ( .A1(n3576), .A2(\vrf/regTable[5][73] ), .B1(n3595), .B2(
        \vrf/regTable[7][73] ), .ZN(n7398) );
  AOI22D1BWP U7197 ( .A1(n8285), .A2(\vrf/regTable[4][73] ), .B1(n3596), .B2(
        \vrf/regTable[6][73] ), .ZN(n7397) );
  AOI22D1BWP U7198 ( .A1(n3579), .A2(\vrf/regTable[1][73] ), .B1(n3599), .B2(
        \vrf/regTable[3][73] ), .ZN(n7396) );
  AOI22D1BWP U7199 ( .A1(n8278), .A2(\vrf/regTable[0][73] ), .B1(n3594), .B2(
        \vrf/regTable[2][73] ), .ZN(n7395) );
  ND4D1BWP U7200 ( .A1(n7971), .A2(n7972), .A3(n7973), .A4(n7974), .ZN(
        vectorData1[217]) );
  AOI22D1BWP U7201 ( .A1(n3576), .A2(\vrf/regTable[5][217] ), .B1(n3595), .B2(
        \vrf/regTable[7][217] ), .ZN(n7974) );
  AOI22D1BWP U7202 ( .A1(n3574), .A2(\vrf/regTable[4][217] ), .B1(n3596), .B2(
        \vrf/regTable[6][217] ), .ZN(n7973) );
  AOI22D1BWP U7203 ( .A1(n3579), .A2(\vrf/regTable[1][217] ), .B1(n3599), .B2(
        \vrf/regTable[3][217] ), .ZN(n7972) );
  AOI22D1BWP U7204 ( .A1(n3581), .A2(\vrf/regTable[0][217] ), .B1(n3594), .B2(
        \vrf/regTable[2][217] ), .ZN(n7971) );
  AOI22D1BWP U7205 ( .A1(n5233), .A2(vectorData1[185]), .B1(n5184), .B2(
        vectorData1[25]), .ZN(n5082) );
  ND4D1BWP U7206 ( .A1(n7203), .A2(n7204), .A3(n7205), .A4(n7206), .ZN(
        vectorData1[25]) );
  AOI22D1BWP U7207 ( .A1(n3576), .A2(\vrf/regTable[5][25] ), .B1(n3595), .B2(
        \vrf/regTable[7][25] ), .ZN(n7206) );
  AOI22D1BWP U7208 ( .A1(n7115), .A2(\vrf/regTable[4][25] ), .B1(n3596), .B2(
        \vrf/regTable[6][25] ), .ZN(n7205) );
  AOI22D1BWP U7209 ( .A1(n3579), .A2(\vrf/regTable[1][25] ), .B1(n3599), .B2(
        \vrf/regTable[3][25] ), .ZN(n7204) );
  AOI22D1BWP U7210 ( .A1(n7108), .A2(\vrf/regTable[0][25] ), .B1(n3594), .B2(
        \vrf/regTable[2][25] ), .ZN(n7203) );
  ND4D1BWP U7211 ( .A1(n7843), .A2(n7844), .A3(n7845), .A4(n7846), .ZN(
        vectorData1[185]) );
  AOI22D1BWP U7212 ( .A1(n3576), .A2(\vrf/regTable[5][185] ), .B1(n3595), .B2(
        \vrf/regTable[7][185] ), .ZN(n7846) );
  AOI22D1BWP U7213 ( .A1(n3574), .A2(\vrf/regTable[4][185] ), .B1(n3596), .B2(
        \vrf/regTable[6][185] ), .ZN(n7845) );
  AOI22D1BWP U7214 ( .A1(n3579), .A2(\vrf/regTable[1][185] ), .B1(n3599), .B2(
        \vrf/regTable[3][185] ), .ZN(n7844) );
  AOI22D1BWP U7215 ( .A1(n3581), .A2(\vrf/regTable[0][185] ), .B1(n3594), .B2(
        \vrf/regTable[2][185] ), .ZN(n7843) );
  AOI22D1BWP U7216 ( .A1(n5213), .A2(vectorData1[105]), .B1(n5230), .B2(
        vectorData1[169]), .ZN(n5083) );
  ND4D1BWP U7217 ( .A1(n7779), .A2(n7780), .A3(n7781), .A4(n7782), .ZN(
        vectorData1[169]) );
  AOI22D1BWP U7218 ( .A1(n3576), .A2(\vrf/regTable[5][169] ), .B1(n3567), .B2(
        \vrf/regTable[7][169] ), .ZN(n7782) );
  AOI22D1BWP U7219 ( .A1(n8285), .A2(\vrf/regTable[4][169] ), .B1(n3570), .B2(
        \vrf/regTable[6][169] ), .ZN(n7781) );
  AOI22D1BWP U7220 ( .A1(n3579), .A2(\vrf/regTable[1][169] ), .B1(n3575), .B2(
        \vrf/regTable[3][169] ), .ZN(n7780) );
  AOI22D1BWP U7221 ( .A1(n8278), .A2(\vrf/regTable[0][169] ), .B1(n3572), .B2(
        \vrf/regTable[2][169] ), .ZN(n7779) );
  ND4D1BWP U7222 ( .A1(n7523), .A2(n7524), .A3(n7525), .A4(n7526), .ZN(
        vectorData1[105]) );
  AOI22D1BWP U7223 ( .A1(n3576), .A2(\vrf/regTable[5][105] ), .B1(n3595), .B2(
        \vrf/regTable[7][105] ), .ZN(n7526) );
  AOI22D1BWP U7224 ( .A1(n3574), .A2(\vrf/regTable[4][105] ), .B1(n3596), .B2(
        \vrf/regTable[6][105] ), .ZN(n7525) );
  AOI22D1BWP U7225 ( .A1(n3579), .A2(\vrf/regTable[1][105] ), .B1(n3575), .B2(
        \vrf/regTable[3][105] ), .ZN(n7524) );
  AOI22D1BWP U7226 ( .A1(n3581), .A2(\vrf/regTable[0][105] ), .B1(n3594), .B2(
        \vrf/regTable[2][105] ), .ZN(n7523) );
  ND4D1BWP U7227 ( .A1(n7715), .A2(n7716), .A3(n7717), .A4(n7718), .ZN(
        vectorData1[153]) );
  AOI22D1BWP U7228 ( .A1(n3576), .A2(\vrf/regTable[5][153] ), .B1(n3595), .B2(
        \vrf/regTable[7][153] ), .ZN(n7718) );
  AOI22D1BWP U7229 ( .A1(n7115), .A2(\vrf/regTable[4][153] ), .B1(n3596), .B2(
        \vrf/regTable[6][153] ), .ZN(n7717) );
  AOI22D1BWP U7230 ( .A1(n3579), .A2(\vrf/regTable[1][153] ), .B1(n3575), .B2(
        \vrf/regTable[3][153] ), .ZN(n7716) );
  AOI22D1BWP U7231 ( .A1(n7108), .A2(\vrf/regTable[0][153] ), .B1(n3594), .B2(
        \vrf/regTable[2][153] ), .ZN(n7715) );
  ND4D1BWP U7232 ( .A1(n7459), .A2(n7460), .A3(n7461), .A4(n7462), .ZN(
        vectorData1[89]) );
  AOI22D1BWP U7233 ( .A1(n7117), .A2(\vrf/regTable[5][89] ), .B1(n3567), .B2(
        \vrf/regTable[7][89] ), .ZN(n7462) );
  AOI22D1BWP U7234 ( .A1(n7115), .A2(\vrf/regTable[4][89] ), .B1(n3570), .B2(
        \vrf/regTable[6][89] ), .ZN(n7461) );
  AOI22D1BWP U7235 ( .A1(n7112), .A2(\vrf/regTable[1][89] ), .B1(n3575), .B2(
        \vrf/regTable[3][89] ), .ZN(n7460) );
  AOI22D1BWP U7236 ( .A1(n7108), .A2(\vrf/regTable[0][89] ), .B1(n3572), .B2(
        \vrf/regTable[2][89] ), .ZN(n7459) );
  ND4D1BWP U7237 ( .A1(n8099), .A2(n8100), .A3(n8101), .A4(n8102), .ZN(
        vectorData1[249]) );
  AOI22D1BWP U7238 ( .A1(n3576), .A2(\vrf/regTable[5][249] ), .B1(n7118), .B2(
        \vrf/regTable[7][249] ), .ZN(n8102) );
  AOI22D1BWP U7239 ( .A1(n3574), .A2(\vrf/regTable[4][249] ), .B1(n7116), .B2(
        \vrf/regTable[6][249] ), .ZN(n8101) );
  AOI22D1BWP U7240 ( .A1(n3579), .A2(\vrf/regTable[1][249] ), .B1(n7114), .B2(
        \vrf/regTable[3][249] ), .ZN(n8100) );
  AOI22D1BWP U7241 ( .A1(n3581), .A2(\vrf/regTable[0][249] ), .B1(n7110), .B2(
        \vrf/regTable[2][249] ), .ZN(n8099) );
  AOI22D1BWP U7242 ( .A1(n3576), .A2(\vrf/regTable[5][57] ), .B1(n3567), .B2(
        \vrf/regTable[7][57] ), .ZN(n7334) );
  AOI22D1BWP U7243 ( .A1(n8285), .A2(\vrf/regTable[4][57] ), .B1(n3570), .B2(
        \vrf/regTable[6][57] ), .ZN(n7333) );
  AOI22D1BWP U7244 ( .A1(n3579), .A2(\vrf/regTable[1][57] ), .B1(n3575), .B2(
        \vrf/regTable[3][57] ), .ZN(n7332) );
  AOI22D1BWP U7245 ( .A1(n8278), .A2(\vrf/regTable[0][57] ), .B1(n3572), .B2(
        \vrf/regTable[2][57] ), .ZN(n7331) );
  AOI22D1BWP U7246 ( .A1(n7117), .A2(\vrf/regTable[5][121] ), .B1(n3567), .B2(
        \vrf/regTable[7][121] ), .ZN(n7590) );
  AOI22D1BWP U7247 ( .A1(n7115), .A2(\vrf/regTable[4][121] ), .B1(n3570), .B2(
        \vrf/regTable[6][121] ), .ZN(n7589) );
  AOI22D1BWP U7248 ( .A1(n7112), .A2(\vrf/regTable[1][121] ), .B1(n3599), .B2(
        \vrf/regTable[3][121] ), .ZN(n7588) );
  AOI22D1BWP U7249 ( .A1(n7108), .A2(\vrf/regTable[0][121] ), .B1(n3572), .B2(
        \vrf/regTable[2][121] ), .ZN(n7587) );
  AO222D1BWP U7250 ( .A1(n4550), .A2(n5495), .B1(n3650), .B2(n5357), .C1(
        vectorToLoad[91]), .C2(n4631), .Z(N4308) );
  NR2XD0BWP U7251 ( .A1(n5290), .A2(\intadd_34/A[0] ), .ZN(n5495) );
  AO222D1BWP U7252 ( .A1(n4550), .A2(n5426), .B1(n3650), .B2(n5308), .C1(
        vectorToLoad[68]), .C2(n3668), .Z(N4285) );
  NR2XD0BWP U7253 ( .A1(n5288), .A2(n4665), .ZN(n5426) );
  AO21D1BWP U7254 ( .A1(nextInstrAddr[6]), .A2(n4061), .B(n3855), .Z(N4140) );
  AOI211XD0BWP U7255 ( .A1(n4661), .A2(n3854), .B(n3903), .C(n3614), .ZN(n3855) );
  IOA21D1BWP U7256 ( .A1(nextInstrAddr[7]), .A2(n4061), .B(n3904), .ZN(N4141)
         );
  OAI211D1BWP U7257 ( .A1(n3903), .A2(result[7]), .B(n4068), .C(n3918), .ZN(
        n3904) );
  AO222D1BWP U7258 ( .A1(n4550), .A2(n5429), .B1(n3650), .B2(n5310), .C1(
        vectorToLoad[69]), .C2(n3669), .Z(N4286) );
  NR2XD0BWP U7259 ( .A1(n5288), .A2(n4664), .ZN(n5429) );
  AO222D1BWP U7260 ( .A1(n4550), .A2(n5432), .B1(n3650), .B2(n5312), .C1(
        vectorToLoad[70]), .C2(n3669), .Z(N4287) );
  NR2XD0BWP U7261 ( .A1(n5288), .A2(n4661), .ZN(n5432) );
  AO21D1BWP U7262 ( .A1(nextInstrAddr[8]), .A2(n4061), .B(n3919), .Z(N4142) );
  AOI211XD0BWP U7263 ( .A1(n4652), .A2(n3918), .B(n4974), .C(n3614), .ZN(n3919) );
  AO222D1BWP U7264 ( .A1(n4550), .A2(n5422), .B1(n5304), .B2(n3650), .C1(
        vectorToLoad[66]), .C2(n3668), .Z(N4283) );
  NR2XD0BWP U7265 ( .A1(n5288), .A2(n4668), .ZN(n5422) );
  AO222D1BWP U7266 ( .A1(n4550), .A2(n5435), .B1(n3650), .B2(n5314), .C1(
        vectorToLoad[71]), .C2(n3668), .Z(N4288) );
  NR2XD0BWP U7267 ( .A1(n5288), .A2(n4655), .ZN(n5435) );
  AO222D1BWP U7268 ( .A1(n4550), .A2(n5438), .B1(n3650), .B2(n5316), .C1(
        vectorToLoad[72]), .C2(n3669), .Z(N4289) );
  NR2XD0BWP U7269 ( .A1(n5288), .A2(n4652), .ZN(n5438) );
  IOA21D1BWP U7270 ( .A1(n4061), .A2(nextInstrAddr[9]), .B(n3926), .ZN(N4143)
         );
  OAI211D1BWP U7271 ( .A1(n4974), .A2(result[9]), .B(n4068), .C(n4975), .ZN(
        n3926) );
  AO222D1BWP U7272 ( .A1(n4550), .A2(n5441), .B1(n3650), .B2(n5318), .C1(
        vectorToLoad[73]), .C2(n3669), .Z(N4290) );
  NR2XD0BWP U7273 ( .A1(n5288), .A2(n4651), .ZN(n5441) );
  AO222D1BWP U7274 ( .A1(n4550), .A2(n5444), .B1(n3650), .B2(n5320), .C1(
        vectorToLoad[74]), .C2(n3668), .Z(N4291) );
  NR2XD0BWP U7275 ( .A1(n5288), .A2(n4699), .ZN(n5444) );
  AO222D1BWP U7276 ( .A1(n4550), .A2(n5420), .B1(n5301), .B2(n3650), .C1(
        vectorToLoad[65]), .C2(n3669), .Z(N4282) );
  NR2XD0BWP U7277 ( .A1(n5288), .A2(n4643), .ZN(n5420) );
  IOA21D1BWP U7278 ( .A1(nextInstrAddr[5]), .A2(n4061), .B(n3845), .ZN(N4139)
         );
  OAI211D1BWP U7279 ( .A1(n4973), .A2(result[5]), .B(n4068), .C(n3854), .ZN(
        n3845) );
  AO222D1BWP U7280 ( .A1(n4550), .A2(n5447), .B1(n3650), .B2(n5322), .C1(
        vectorToLoad[75]), .C2(n3668), .Z(N4292) );
  NR2XD0BWP U7281 ( .A1(n5288), .A2(\intadd_34/A[0] ), .ZN(n5447) );
  OAI22D1BWP U7282 ( .A1(n4977), .A2(n3614), .B1(n4064), .B2(n3861), .ZN(N4145) );
  AOI32D1BWP U7283 ( .A1(result[10]), .A2(n4978), .A3(n4976), .B1(result[11]), 
        .B2(n4978), .ZN(n4977) );
  AO222D1BWP U7284 ( .A1(n4550), .A2(n5450), .B1(n3650), .B2(n5324), .C1(
        vectorToLoad[76]), .C2(n3668), .Z(N4293) );
  NR2XD0BWP U7285 ( .A1(n5288), .A2(\intadd_34/A[1] ), .ZN(n5450) );
  NR2XD0BWP U7286 ( .A1(n5286), .A2(n5285), .ZN(n5414) );
  AO222D1BWP U7287 ( .A1(n4550), .A2(n5453), .B1(n3650), .B2(n5326), .C1(
        vectorToLoad[77]), .C2(n3669), .Z(N4294) );
  NR2XD0BWP U7288 ( .A1(n5288), .A2(\intadd_34/A[2] ), .ZN(n5453) );
  AOI22D1BWP U7289 ( .A1(result[12]), .A2(n4978), .B1(n4981), .B2(
        \intadd_34/A[1] ), .ZN(n4979) );
  AO222D1BWP U7290 ( .A1(n4550), .A2(n5456), .B1(n3650), .B2(n5328), .C1(
        vectorToLoad[78]), .C2(n3668), .Z(N4295) );
  NR2XD0BWP U7291 ( .A1(n5288), .A2(\intadd_34/A[3] ), .ZN(n5456) );
  AO222D1BWP U7292 ( .A1(n4550), .A2(n5459), .B1(n3650), .B2(n5330), .C1(
        vectorToLoad[79]), .C2(n3669), .Z(N4296) );
  NR2XD0BWP U7293 ( .A1(n5288), .A2(n6037), .ZN(n5459) );
  OAI22D1BWP U7294 ( .A1(n4982), .A2(n3614), .B1(n4064), .B2(n4063), .ZN(N4147) );
  AOI32D1BWP U7295 ( .A1(result[12]), .A2(n4983), .A3(n4981), .B1(result[13]), 
        .B2(n4983), .ZN(n4982) );
  AO222D1BWP U7296 ( .A1(n3668), .A2(vectorToLoad[80]), .B1(n5462), .B2(n3667), 
        .C1(n5289), .C2(n3650), .Z(N4297) );
  AO222D1BWP U7297 ( .A1(n3669), .A2(vectorToLoad[63]), .B1(n5412), .B2(n3649), 
        .C1(n4549), .C2(n5553), .Z(N4280) );
  OAI31D1BWP U7298 ( .A1(n4984), .A2(n4069), .A3(n3614), .B(n4989), .ZN(N4148)
         );
  NR2XD0BWP U7299 ( .A1(n4067), .A2(result[14]), .ZN(n4069) );
  AO222D1BWP U7300 ( .A1(n4550), .A2(n5465), .B1(n3650), .B2(n5387), .C1(
        vectorToLoad[81]), .C2(n3668), .Z(N4298) );
  NR2XD0BWP U7301 ( .A1(n5290), .A2(n4643), .ZN(n5465) );
  AO222D1BWP U7302 ( .A1(n4550), .A2(n5468), .B1(n3650), .B2(n5389), .C1(
        vectorToLoad[82]), .C2(n4631), .Z(N4299) );
  NR2XD0BWP U7303 ( .A1(n5290), .A2(n4668), .ZN(n5468) );
  OAI21D1BWP U7304 ( .A1(n4985), .A2(n3614), .B(n4391), .ZN(N4149) );
  NR2XD0BWP U7305 ( .A1(\intadd_34/A[3] ), .A2(n4983), .ZN(n4984) );
  ND3D1BWP U7306 ( .A1(result[11]), .A2(result[10]), .A3(n4976), .ZN(n4978) );
  NR2XD0BWP U7307 ( .A1(n3918), .A2(n4652), .ZN(n4974) );
  NR2XD0BWP U7308 ( .A1(n3854), .A2(n4661), .ZN(n3903) );
  MAOI222D1BWP U7309 ( .A(n4969), .B(cycles[3]), .C(result[3]), .ZN(n4971) );
  AO222D1BWP U7310 ( .A1(n4550), .A2(n5471), .B1(n3650), .B2(n5391), .C1(
        vectorToLoad[83]), .C2(n4631), .Z(N4300) );
  NR2XD0BWP U7311 ( .A1(n5290), .A2(n6011), .ZN(n5471) );
  AO222D1BWP U7312 ( .A1(n3669), .A2(vectorToLoad[62]), .B1(n5410), .B2(n3649), 
        .C1(n4549), .C2(n5552), .Z(N4279) );
  AO222D1BWP U7313 ( .A1(n4550), .A2(n5474), .B1(n3650), .B2(n5341), .C1(
        vectorToLoad[84]), .C2(n4631), .Z(N4301) );
  NR2XD0BWP U7314 ( .A1(n5290), .A2(n4665), .ZN(n5474) );
  AO222D1BWP U7315 ( .A1(n4550), .A2(n5477), .B1(n3650), .B2(n5394), .C1(
        vectorToLoad[85]), .C2(n4631), .Z(N4302) );
  NR2XD0BWP U7316 ( .A1(n5290), .A2(n4664), .ZN(n5477) );
  AO222D1BWP U7317 ( .A1(n3669), .A2(vectorToLoad[61]), .B1(n5408), .B2(n3649), 
        .C1(n4549), .C2(n5551), .Z(N4278) );
  AO222D1BWP U7318 ( .A1(n4550), .A2(n5480), .B1(n3650), .B2(n5396), .C1(
        vectorToLoad[86]), .C2(n4631), .Z(N4303) );
  NR2XD0BWP U7319 ( .A1(n5290), .A2(n4661), .ZN(n5480) );
  AO222D1BWP U7320 ( .A1(n4550), .A2(n5483), .B1(n3650), .B2(n5398), .C1(
        vectorToLoad[87]), .C2(n4631), .Z(N4304) );
  NR2XD0BWP U7321 ( .A1(n5290), .A2(n4655), .ZN(n5483) );
  AO222D1BWP U7322 ( .A1(n4550), .A2(n5486), .B1(n3650), .B2(n5400), .C1(
        vectorToLoad[88]), .C2(n4631), .Z(N4305) );
  NR2XD0BWP U7323 ( .A1(n5290), .A2(n4652), .ZN(n5486) );
  AO222D1BWP U7324 ( .A1(n3668), .A2(vectorToLoad[60]), .B1(n5406), .B2(n3649), 
        .C1(n4549), .C2(n5550), .Z(N4277) );
  ND4D1BWP U7325 ( .A1(n5212), .A2(n5211), .A3(n5210), .A4(n5209), .ZN(N4204)
         );
  AOI31D1BWP U7326 ( .A1(n5204), .A2(n5206), .A3(n5205), .B(n3661), .ZN(n5207)
         );
  AOI22D1BWP U7327 ( .A1(vectorData2[220]), .A2(n5228), .B1(vectorData2[156]), 
        .B2(n5232), .ZN(n5205) );
  AOI22D1BWP U7328 ( .A1(vectorData2[140]), .A2(n5226), .B1(vectorData2[44]), 
        .B2(n3601), .ZN(n5206) );
  OA211D1BWP U7329 ( .A1(n5203), .A2(n3674), .B(n5202), .C(n5201), .Z(n5204)
         );
  AOI22D1BWP U7330 ( .A1(vectorData2[204]), .A2(n5227), .B1(vectorData2[172]), 
        .B2(n5230), .ZN(n5201) );
  AOI22D1BWP U7331 ( .A1(vectorData2[252]), .A2(n5229), .B1(vectorData2[188]), 
        .B2(n5233), .ZN(n5202) );
  AOI22D1BWP U7332 ( .A1(vectorData2[92]), .A2(n4684), .B1(vectorData2[12]), 
        .B2(n4681), .ZN(n5208) );
  AOI22D1BWP U7333 ( .A1(vectorData2[108]), .A2(n4683), .B1(vectorData2[28]), 
        .B2(n4685), .ZN(n5210) );
  AOI22D1BWP U7334 ( .A1(vectorData2[76]), .A2(n4682), .B1(scalarData2[12]), 
        .B2(n4688), .ZN(n5211) );
  AOI22D1BWP U7335 ( .A1(vectorData2[236]), .A2(n4694), .B1(vectorData2[60]), 
        .B2(n4686), .ZN(n5212) );
  AO222D1BWP U7336 ( .A1(n4550), .A2(n5489), .B1(n3650), .B2(n5352), .C1(
        vectorToLoad[89]), .C2(n4631), .Z(N4306) );
  NR2XD0BWP U7337 ( .A1(n5290), .A2(n4651), .ZN(n5489) );
  AO222D1BWP U7338 ( .A1(n4550), .A2(n5492), .B1(n3650), .B2(n5403), .C1(
        vectorToLoad[90]), .C2(n4631), .Z(N4307) );
  NR2XD0BWP U7339 ( .A1(n5290), .A2(n4699), .ZN(n5492) );
  AO222D1BWP U7340 ( .A1(n4550), .A2(n5424), .B1(n5306), .B2(n3650), .C1(
        vectorToLoad[67]), .C2(n3669), .Z(N4284) );
  NR2XD0BWP U7341 ( .A1(n5288), .A2(n6011), .ZN(n5424) );
  AO222D1BWP U7342 ( .A1(n3668), .A2(vectorToLoad[44]), .B1(n4549), .B2(n5532), 
        .C1(n3649), .C2(n5324), .Z(N4261) );
  OAI211D1BWP U7343 ( .A1(n5437), .A2(n4407), .B(n5377), .C(n4535), .ZN(N4385)
         );
  AOI22D1BWP U7344 ( .A1(n3669), .A2(vectorToLoad[167]), .B1(n5415), .B2(n5527), .ZN(n5377) );
  OAI211D1BWP U7345 ( .A1(n5440), .A2(n4407), .B(n5378), .C(n4535), .ZN(N4386)
         );
  AOI22D1BWP U7346 ( .A1(n3668), .A2(vectorToLoad[168]), .B1(n5415), .B2(n5528), .ZN(n5378) );
  AO222D1BWP U7347 ( .A1(n3644), .A2(n4548), .B1(n5530), .B2(n4628), .C1(n3669), .C2(vectorToLoad[106]), .Z(N4323) );
  OAI211D1BWP U7348 ( .A1(n5443), .A2(n4407), .B(n5379), .C(n4535), .ZN(N4387)
         );
  AOI22D1BWP U7349 ( .A1(n3669), .A2(vectorToLoad[169]), .B1(n5415), .B2(n5529), .ZN(n5379) );
  AO222D1BWP U7350 ( .A1(n3668), .A2(vectorToLoad[43]), .B1(n4549), .B2(n5531), 
        .C1(n3649), .C2(n5322), .Z(N4260) );
  OAI211D1BWP U7351 ( .A1(n5446), .A2(n4407), .B(n5380), .C(n4535), .ZN(N4388)
         );
  AOI22D1BWP U7352 ( .A1(n3668), .A2(vectorToLoad[170]), .B1(n5415), .B2(n5530), .ZN(n5380) );
  OAI211D1BWP U7353 ( .A1(n5449), .A2(n4407), .B(n5381), .C(n4535), .ZN(N4389)
         );
  AOI22D1BWP U7354 ( .A1(n3669), .A2(vectorToLoad[171]), .B1(n5415), .B2(n5531), .ZN(n5381) );
  OAI211D1BWP U7355 ( .A1(n5452), .A2(n4407), .B(n5382), .C(n4535), .ZN(N4390)
         );
  AOI22D1BWP U7356 ( .A1(n3668), .A2(vectorToLoad[172]), .B1(n5415), .B2(n5532), .ZN(n5382) );
  AO222D1BWP U7357 ( .A1(n3669), .A2(vectorToLoad[42]), .B1(n4549), .B2(n5530), 
        .C1(n3649), .C2(n5320), .Z(N4259) );
  NR2XD0BWP U7358 ( .A1(n4699), .A2(n5282), .ZN(n5530) );
  OAI211D1BWP U7359 ( .A1(n5455), .A2(n4407), .B(n5383), .C(n4535), .ZN(N4391)
         );
  AOI22D1BWP U7360 ( .A1(n3668), .A2(vectorToLoad[173]), .B1(n5415), .B2(n5533), .ZN(n5383) );
  AO222D1BWP U7361 ( .A1(n3645), .A2(n4548), .B1(n5531), .B2(n3667), .C1(n4631), .C2(vectorToLoad[107]), .Z(N4324) );
  NR2XD0BWP U7362 ( .A1(\intadd_34/A[0] ), .A2(n5282), .ZN(n5531) );
  OAI211D1BWP U7363 ( .A1(n5458), .A2(n4407), .B(n5384), .C(n4535), .ZN(N4392)
         );
  AOI22D1BWP U7364 ( .A1(n3668), .A2(vectorToLoad[174]), .B1(n5415), .B2(n5534), .ZN(n5384) );
  OAI211D1BWP U7365 ( .A1(n5461), .A2(n4407), .B(n5385), .C(n4535), .ZN(N4393)
         );
  AOI22D1BWP U7366 ( .A1(n3668), .A2(vectorToLoad[175]), .B1(n5415), .B2(n5535), .ZN(n5385) );
  OAI211D1BWP U7367 ( .A1(n5464), .A2(n4407), .B(n5386), .C(n4535), .ZN(N4394)
         );
  AOI22D1BWP U7368 ( .A1(vectorToLoad[176]), .A2(n3668), .B1(n5415), .B2(n5536), .ZN(n5386) );
  AO222D1BWP U7369 ( .A1(n3668), .A2(vectorToLoad[41]), .B1(n4549), .B2(n5529), 
        .C1(n3649), .C2(n5318), .Z(N4258) );
  OAI211D1BWP U7370 ( .A1(n5467), .A2(n4407), .B(n5388), .C(n4535), .ZN(N4395)
         );
  AOI22D1BWP U7371 ( .A1(n3668), .A2(vectorToLoad[177]), .B1(n5415), .B2(n5539), .ZN(n5388) );
  OAI211D1BWP U7372 ( .A1(n5470), .A2(n4407), .B(n5390), .C(n4535), .ZN(N4396)
         );
  AOI22D1BWP U7373 ( .A1(n3668), .A2(vectorToLoad[178]), .B1(n5415), .B2(n5540), .ZN(n5390) );
  AO222D1BWP U7374 ( .A1(n3646), .A2(n4548), .B1(n5532), .B2(n4628), .C1(n3668), .C2(vectorToLoad[108]), .Z(N4325) );
  NR2XD0BWP U7375 ( .A1(\intadd_34/A[1] ), .A2(n5282), .ZN(n5532) );
  NR2XD0BWP U7376 ( .A1(n3679), .A2(n5279), .ZN(n5324) );
  OAI211D1BWP U7377 ( .A1(n5473), .A2(n4407), .B(n5392), .C(n4535), .ZN(N4397)
         );
  AOI22D1BWP U7378 ( .A1(n3668), .A2(vectorToLoad[179]), .B1(n5415), .B2(n5541), .ZN(n5392) );
  AO222D1BWP U7379 ( .A1(n3668), .A2(vectorToLoad[40]), .B1(n4549), .B2(n5528), 
        .C1(n3649), .C2(n5316), .Z(N4257) );
  OAI211D1BWP U7380 ( .A1(n5476), .A2(n4407), .B(n5393), .C(n4535), .ZN(N4398)
         );
  AOI22D1BWP U7381 ( .A1(n3668), .A2(vectorToLoad[180]), .B1(n5415), .B2(n5542), .ZN(n5393) );
  OAI211D1BWP U7382 ( .A1(n5479), .A2(n4407), .B(n5395), .C(n4535), .ZN(N4399)
         );
  AOI22D1BWP U7383 ( .A1(n3668), .A2(vectorToLoad[181]), .B1(n5415), .B2(n5543), .ZN(n5395) );
  OAI211D1BWP U7384 ( .A1(n5482), .A2(n4407), .B(n5397), .C(n4535), .ZN(N4400)
         );
  AOI22D1BWP U7385 ( .A1(n3668), .A2(vectorToLoad[182]), .B1(n5415), .B2(n5544), .ZN(n5397) );
  AO222D1BWP U7386 ( .A1(n3669), .A2(vectorToLoad[39]), .B1(n4549), .B2(n5527), 
        .C1(n3649), .C2(n5314), .Z(N4256) );
  OAI211D1BWP U7387 ( .A1(n5485), .A2(n4407), .B(n5399), .C(n4535), .ZN(N4401)
         );
  AOI22D1BWP U7388 ( .A1(n3668), .A2(vectorToLoad[183]), .B1(n5415), .B2(n5545), .ZN(n5399) );
  OAI211D1BWP U7389 ( .A1(n5488), .A2(n4407), .B(n5401), .C(n4535), .ZN(N4402)
         );
  AOI22D1BWP U7390 ( .A1(n3668), .A2(vectorToLoad[184]), .B1(n5415), .B2(n5546), .ZN(n5401) );
  AO222D1BWP U7391 ( .A1(n3647), .A2(n4548), .B1(n5533), .B2(n3667), .C1(n3668), .C2(vectorToLoad[109]), .Z(N4326) );
  OAI211D1BWP U7392 ( .A1(n5491), .A2(n4407), .B(n5402), .C(n4535), .ZN(N4403)
         );
  AOI22D1BWP U7393 ( .A1(n3668), .A2(vectorToLoad[185]), .B1(n5415), .B2(n5547), .ZN(n5402) );
  AO222D1BWP U7394 ( .A1(n3669), .A2(vectorToLoad[38]), .B1(n4549), .B2(n5526), 
        .C1(n3649), .C2(n5312), .Z(N4255) );
  OAI211D1BWP U7395 ( .A1(n5494), .A2(n4407), .B(n5404), .C(n4535), .ZN(N4404)
         );
  AOI22D1BWP U7396 ( .A1(n3668), .A2(vectorToLoad[186]), .B1(n5415), .B2(n5548), .ZN(n5404) );
  OAI211D1BWP U7397 ( .A1(n5497), .A2(n4407), .B(n5405), .C(n4535), .ZN(N4405)
         );
  AOI22D1BWP U7398 ( .A1(n3668), .A2(vectorToLoad[187]), .B1(n5415), .B2(n5549), .ZN(n5405) );
  OAI211D1BWP U7399 ( .A1(n5500), .A2(n4407), .B(n5407), .C(n4535), .ZN(N4406)
         );
  AOI22D1BWP U7400 ( .A1(n3668), .A2(vectorToLoad[188]), .B1(n5415), .B2(n5550), .ZN(n5407) );
  AO222D1BWP U7401 ( .A1(n3668), .A2(vectorToLoad[37]), .B1(n4549), .B2(n5525), 
        .C1(n3649), .C2(n5310), .Z(N4254) );
  OAI211D1BWP U7402 ( .A1(n5434), .A2(n4407), .B(n5376), .C(n4535), .ZN(N4384)
         );
  AOI22D1BWP U7403 ( .A1(n3668), .A2(vectorToLoad[166]), .B1(n5415), .B2(n5526), .ZN(n5376) );
  OAI211D1BWP U7404 ( .A1(n5461), .A2(n4405), .B(n5332), .C(n4535), .ZN(N4361)
         );
  AOI22D1BWP U7405 ( .A1(result[15]), .A2(n5331), .B1(n3668), .B2(
        vectorToLoad[143]), .ZN(n5332) );
  NR2XD0BWP U7406 ( .A1(n5302), .A2(n5509), .ZN(n5331) );
  OAI211D1BWP U7407 ( .A1(n5464), .A2(n4405), .B(n5333), .C(n4535), .ZN(N4362)
         );
  AOI22D1BWP U7408 ( .A1(n3669), .A2(vectorToLoad[144]), .B1(n5415), .B2(n5462), .ZN(n5333) );
  NR2XD0BWP U7409 ( .A1(cycles[1]), .A2(n5284), .ZN(n5462) );
  AO211D1BWP U7410 ( .A1(n4073), .A2(scalarData1[8]), .B(n3921), .C(n3920), 
        .Z(N4184) );
  AO22D1BWP U7411 ( .A1(n4072), .A2(vectorData1[8]), .B1(n4071), .B2(Addr[8]), 
        .Z(n3920) );
  ND4D1BWP U7412 ( .A1(n7151), .A2(n7152), .A3(n7153), .A4(n7154), .ZN(
        vectorData1[8]) );
  AOI22D1BWP U7413 ( .A1(n3576), .A2(\vrf/regTable[5][8] ), .B1(n3595), .B2(
        \vrf/regTable[7][8] ), .ZN(n7154) );
  AOI22D1BWP U7414 ( .A1(n3574), .A2(\vrf/regTable[4][8] ), .B1(n3596), .B2(
        \vrf/regTable[6][8] ), .ZN(n7153) );
  AOI22D1BWP U7415 ( .A1(n3579), .A2(\vrf/regTable[1][8] ), .B1(n3599), .B2(
        \vrf/regTable[3][8] ), .ZN(n7152) );
  AOI22D1BWP U7416 ( .A1(n3581), .A2(\vrf/regTable[0][8] ), .B1(n3594), .B2(
        \vrf/regTable[2][8] ), .ZN(n7151) );
  AOI31D1BWP U7417 ( .A1(n5078), .A2(n5077), .A3(n5079), .B(n4070), .ZN(n3921)
         );
  AOI22D1BWP U7418 ( .A1(n5233), .A2(vectorData1[184]), .B1(n3601), .B2(
        vectorData1[40]), .ZN(n5079) );
  ND4D1BWP U7419 ( .A1(n7263), .A2(n7264), .A3(n7265), .A4(n7266), .ZN(
        vectorData1[40]) );
  AOI22D1BWP U7420 ( .A1(n3576), .A2(\vrf/regTable[5][40] ), .B1(n3595), .B2(
        \vrf/regTable[7][40] ), .ZN(n7266) );
  AOI22D1BWP U7421 ( .A1(n3574), .A2(\vrf/regTable[4][40] ), .B1(n3596), .B2(
        \vrf/regTable[6][40] ), .ZN(n7265) );
  AOI22D1BWP U7422 ( .A1(n3579), .A2(\vrf/regTable[1][40] ), .B1(n3599), .B2(
        \vrf/regTable[3][40] ), .ZN(n7264) );
  AOI22D1BWP U7423 ( .A1(n3581), .A2(\vrf/regTable[0][40] ), .B1(n3594), .B2(
        \vrf/regTable[2][40] ), .ZN(n7263) );
  ND4D1BWP U7424 ( .A1(n7839), .A2(n7840), .A3(n7841), .A4(n7842), .ZN(
        vectorData1[184]) );
  AOI22D1BWP U7425 ( .A1(n3576), .A2(\vrf/regTable[5][184] ), .B1(n7118), .B2(
        \vrf/regTable[7][184] ), .ZN(n7842) );
  AOI22D1BWP U7426 ( .A1(n3574), .A2(\vrf/regTable[4][184] ), .B1(n7116), .B2(
        \vrf/regTable[6][184] ), .ZN(n7841) );
  AOI22D1BWP U7427 ( .A1(n3579), .A2(\vrf/regTable[1][184] ), .B1(n7114), .B2(
        \vrf/regTable[3][184] ), .ZN(n7840) );
  AOI22D1BWP U7428 ( .A1(n3581), .A2(\vrf/regTable[0][184] ), .B1(n7110), .B2(
        \vrf/regTable[2][184] ), .ZN(n7839) );
  AOI211XD0BWP U7429 ( .A1(n5228), .A2(vectorData1[216]), .B(n5076), .C(n5075), 
        .ZN(n5077) );
  ND4D1BWP U7430 ( .A1(n5074), .A2(n5073), .A3(n5072), .A4(n5071), .ZN(n5075)
         );
  AOI22D1BWP U7431 ( .A1(n5184), .A2(vectorData1[24]), .B1(n5227), .B2(
        vectorData1[200]), .ZN(n5071) );
  ND4D1BWP U7432 ( .A1(n7903), .A2(n7904), .A3(n7905), .A4(n7906), .ZN(
        vectorData1[200]) );
  AOI22D1BWP U7433 ( .A1(n3576), .A2(\vrf/regTable[5][200] ), .B1(n7118), .B2(
        \vrf/regTable[7][200] ), .ZN(n7906) );
  AOI22D1BWP U7434 ( .A1(n3574), .A2(\vrf/regTable[4][200] ), .B1(n7116), .B2(
        \vrf/regTable[6][200] ), .ZN(n7905) );
  AOI22D1BWP U7435 ( .A1(n3579), .A2(\vrf/regTable[1][200] ), .B1(n7114), .B2(
        \vrf/regTable[3][200] ), .ZN(n7904) );
  AOI22D1BWP U7436 ( .A1(n3581), .A2(\vrf/regTable[0][200] ), .B1(n7110), .B2(
        \vrf/regTable[2][200] ), .ZN(n7903) );
  ND4D1BWP U7437 ( .A1(n7199), .A2(n7200), .A3(n7201), .A4(n7202), .ZN(
        vectorData1[24]) );
  AOI22D1BWP U7438 ( .A1(n3576), .A2(\vrf/regTable[5][24] ), .B1(n3567), .B2(
        \vrf/regTable[7][24] ), .ZN(n7202) );
  AOI22D1BWP U7439 ( .A1(n7115), .A2(\vrf/regTable[4][24] ), .B1(n3570), .B2(
        \vrf/regTable[6][24] ), .ZN(n7201) );
  AOI22D1BWP U7440 ( .A1(n3579), .A2(\vrf/regTable[1][24] ), .B1(n3575), .B2(
        \vrf/regTable[3][24] ), .ZN(n7200) );
  AOI22D1BWP U7441 ( .A1(n7108), .A2(\vrf/regTable[0][24] ), .B1(n3572), .B2(
        \vrf/regTable[2][24] ), .ZN(n7199) );
  AOI22D1BWP U7442 ( .A1(n5187), .A2(vectorData1[232]), .B1(n5230), .B2(
        vectorData1[168]), .ZN(n5072) );
  ND4D1BWP U7443 ( .A1(n7775), .A2(n7776), .A3(n7777), .A4(n7778), .ZN(
        vectorData1[168]) );
  AOI22D1BWP U7444 ( .A1(n3576), .A2(\vrf/regTable[5][168] ), .B1(n3595), .B2(
        \vrf/regTable[7][168] ), .ZN(n7778) );
  AOI22D1BWP U7445 ( .A1(n3574), .A2(\vrf/regTable[4][168] ), .B1(n3596), .B2(
        \vrf/regTable[6][168] ), .ZN(n7777) );
  AOI22D1BWP U7446 ( .A1(n3579), .A2(\vrf/regTable[1][168] ), .B1(n3575), .B2(
        \vrf/regTable[3][168] ), .ZN(n7776) );
  AOI22D1BWP U7447 ( .A1(n3581), .A2(\vrf/regTable[0][168] ), .B1(n3594), .B2(
        \vrf/regTable[2][168] ), .ZN(n7775) );
  ND4D1BWP U7448 ( .A1(n8031), .A2(n8032), .A3(n8033), .A4(n8034), .ZN(
        vectorData1[232]) );
  AOI22D1BWP U7449 ( .A1(n3576), .A2(\vrf/regTable[5][232] ), .B1(n3595), .B2(
        \vrf/regTable[7][232] ), .ZN(n8034) );
  AOI22D1BWP U7450 ( .A1(n8285), .A2(\vrf/regTable[4][232] ), .B1(n3596), .B2(
        \vrf/regTable[6][232] ), .ZN(n8033) );
  AOI22D1BWP U7451 ( .A1(n3579), .A2(\vrf/regTable[1][232] ), .B1(n3599), .B2(
        \vrf/regTable[3][232] ), .ZN(n8032) );
  AOI22D1BWP U7452 ( .A1(n8278), .A2(\vrf/regTable[0][232] ), .B1(n3594), .B2(
        \vrf/regTable[2][232] ), .ZN(n8031) );
  AOI22D1BWP U7453 ( .A1(n5226), .A2(vectorData1[136]), .B1(n5229), .B2(
        vectorData1[248]), .ZN(n5073) );
  ND4D1BWP U7454 ( .A1(n8095), .A2(n8096), .A3(n8097), .A4(n8098), .ZN(
        vectorData1[248]) );
  AOI22D1BWP U7455 ( .A1(n3576), .A2(\vrf/regTable[5][248] ), .B1(n3595), .B2(
        \vrf/regTable[7][248] ), .ZN(n8098) );
  AOI22D1BWP U7456 ( .A1(n3574), .A2(\vrf/regTable[4][248] ), .B1(n3596), .B2(
        \vrf/regTable[6][248] ), .ZN(n8097) );
  AOI22D1BWP U7457 ( .A1(n3579), .A2(\vrf/regTable[1][248] ), .B1(n3599), .B2(
        \vrf/regTable[3][248] ), .ZN(n8096) );
  AOI22D1BWP U7458 ( .A1(n3581), .A2(\vrf/regTable[0][248] ), .B1(n3594), .B2(
        \vrf/regTable[2][248] ), .ZN(n8095) );
  ND4D1BWP U7459 ( .A1(n7647), .A2(n7648), .A3(n7649), .A4(n7650), .ZN(
        vectorData1[136]) );
  AOI22D1BWP U7460 ( .A1(n3576), .A2(\vrf/regTable[5][136] ), .B1(n3567), .B2(
        \vrf/regTable[7][136] ), .ZN(n7650) );
  AOI22D1BWP U7461 ( .A1(n3574), .A2(\vrf/regTable[4][136] ), .B1(n3570), .B2(
        \vrf/regTable[6][136] ), .ZN(n7649) );
  AOI22D1BWP U7462 ( .A1(n3579), .A2(\vrf/regTable[1][136] ), .B1(n3599), .B2(
        \vrf/regTable[3][136] ), .ZN(n7648) );
  AOI22D1BWP U7463 ( .A1(n3581), .A2(\vrf/regTable[0][136] ), .B1(n3572), .B2(
        \vrf/regTable[2][136] ), .ZN(n7647) );
  AOI22D1BWP U7464 ( .A1(n5231), .A2(vectorData1[120]), .B1(n5188), .B2(
        vectorData1[56]), .ZN(n5074) );
  ND4D1BWP U7465 ( .A1(n7327), .A2(n7328), .A3(n7329), .A4(n7330), .ZN(
        vectorData1[56]) );
  AOI22D1BWP U7466 ( .A1(n3576), .A2(\vrf/regTable[5][56] ), .B1(n3567), .B2(
        \vrf/regTable[7][56] ), .ZN(n7330) );
  AOI22D1BWP U7467 ( .A1(n3574), .A2(\vrf/regTable[4][56] ), .B1(n3570), .B2(
        \vrf/regTable[6][56] ), .ZN(n7329) );
  AOI22D1BWP U7468 ( .A1(n3579), .A2(\vrf/regTable[1][56] ), .B1(n3575), .B2(
        \vrf/regTable[3][56] ), .ZN(n7328) );
  AOI22D1BWP U7469 ( .A1(n3581), .A2(\vrf/regTable[0][56] ), .B1(n3572), .B2(
        \vrf/regTable[2][56] ), .ZN(n7327) );
  ND4D1BWP U7470 ( .A1(n7583), .A2(n7584), .A3(n7585), .A4(n7586), .ZN(
        vectorData1[120]) );
  AOI22D1BWP U7471 ( .A1(n3576), .A2(\vrf/regTable[5][120] ), .B1(n3595), .B2(
        \vrf/regTable[7][120] ), .ZN(n7586) );
  AOI22D1BWP U7472 ( .A1(n3574), .A2(\vrf/regTable[4][120] ), .B1(n3596), .B2(
        \vrf/regTable[6][120] ), .ZN(n7585) );
  AOI22D1BWP U7473 ( .A1(n3579), .A2(\vrf/regTable[1][120] ), .B1(n3575), .B2(
        \vrf/regTable[3][120] ), .ZN(n7584) );
  AOI22D1BWP U7474 ( .A1(n3581), .A2(\vrf/regTable[0][120] ), .B1(n3594), .B2(
        \vrf/regTable[2][120] ), .ZN(n7583) );
  AO22D1BWP U7475 ( .A1(n5185), .A2(vectorData1[88]), .B1(n5186), .B2(
        vectorData1[72]), .Z(n5076) );
  ND4D1BWP U7476 ( .A1(n7391), .A2(n7392), .A3(n7393), .A4(n7394), .ZN(
        vectorData1[72]) );
  AOI22D1BWP U7477 ( .A1(n3576), .A2(\vrf/regTable[5][72] ), .B1(n3595), .B2(
        \vrf/regTable[7][72] ), .ZN(n7394) );
  AOI22D1BWP U7478 ( .A1(n3574), .A2(\vrf/regTable[4][72] ), .B1(n3596), .B2(
        \vrf/regTable[6][72] ), .ZN(n7393) );
  AOI22D1BWP U7479 ( .A1(n3579), .A2(\vrf/regTable[1][72] ), .B1(n3599), .B2(
        \vrf/regTable[3][72] ), .ZN(n7392) );
  AOI22D1BWP U7480 ( .A1(n3581), .A2(\vrf/regTable[0][72] ), .B1(n3594), .B2(
        \vrf/regTable[2][72] ), .ZN(n7391) );
  ND4D1BWP U7481 ( .A1(n7455), .A2(n7456), .A3(n7457), .A4(n7458), .ZN(
        vectorData1[88]) );
  AOI22D1BWP U7482 ( .A1(n7117), .A2(\vrf/regTable[5][88] ), .B1(n3567), .B2(
        \vrf/regTable[7][88] ), .ZN(n7458) );
  AOI22D1BWP U7483 ( .A1(n7115), .A2(\vrf/regTable[4][88] ), .B1(n3570), .B2(
        \vrf/regTable[6][88] ), .ZN(n7457) );
  AOI22D1BWP U7484 ( .A1(n7112), .A2(\vrf/regTable[1][88] ), .B1(n3575), .B2(
        \vrf/regTable[3][88] ), .ZN(n7456) );
  AOI22D1BWP U7485 ( .A1(n7108), .A2(\vrf/regTable[0][88] ), .B1(n3572), .B2(
        \vrf/regTable[2][88] ), .ZN(n7455) );
  ND4D1BWP U7486 ( .A1(n7967), .A2(n7968), .A3(n7969), .A4(n7970), .ZN(
        vectorData1[216]) );
  AOI22D1BWP U7487 ( .A1(n3576), .A2(\vrf/regTable[5][216] ), .B1(n3595), .B2(
        \vrf/regTable[7][216] ), .ZN(n7970) );
  AOI22D1BWP U7488 ( .A1(n3574), .A2(\vrf/regTable[4][216] ), .B1(n3596), .B2(
        \vrf/regTable[6][216] ), .ZN(n7969) );
  AOI22D1BWP U7489 ( .A1(n3579), .A2(\vrf/regTable[1][216] ), .B1(n3599), .B2(
        \vrf/regTable[3][216] ), .ZN(n7968) );
  AOI22D1BWP U7490 ( .A1(n3581), .A2(\vrf/regTable[0][216] ), .B1(n3594), .B2(
        \vrf/regTable[2][216] ), .ZN(n7967) );
  AOI22D1BWP U7491 ( .A1(n5213), .A2(vectorData1[104]), .B1(n5232), .B2(
        vectorData1[152]), .ZN(n5078) );
  ND4D1BWP U7492 ( .A1(n7711), .A2(n7712), .A3(n7713), .A4(n7714), .ZN(
        vectorData1[152]) );
  AOI22D1BWP U7493 ( .A1(n3576), .A2(\vrf/regTable[5][152] ), .B1(n3595), .B2(
        \vrf/regTable[7][152] ), .ZN(n7714) );
  AOI22D1BWP U7494 ( .A1(n3574), .A2(\vrf/regTable[4][152] ), .B1(n3596), .B2(
        \vrf/regTable[6][152] ), .ZN(n7713) );
  AOI22D1BWP U7495 ( .A1(n3579), .A2(\vrf/regTable[1][152] ), .B1(n3599), .B2(
        \vrf/regTable[3][152] ), .ZN(n7712) );
  AOI22D1BWP U7496 ( .A1(n3581), .A2(\vrf/regTable[0][152] ), .B1(n3594), .B2(
        \vrf/regTable[2][152] ), .ZN(n7711) );
  ND4D1BWP U7497 ( .A1(n7519), .A2(n7520), .A3(n7521), .A4(n7522), .ZN(
        vectorData1[104]) );
  AOI22D1BWP U7498 ( .A1(n3576), .A2(\vrf/regTable[5][104] ), .B1(n3595), .B2(
        \vrf/regTable[7][104] ), .ZN(n7522) );
  AOI22D1BWP U7499 ( .A1(n3574), .A2(\vrf/regTable[4][104] ), .B1(n3596), .B2(
        \vrf/regTable[6][104] ), .ZN(n7521) );
  AOI22D1BWP U7500 ( .A1(n3579), .A2(\vrf/regTable[1][104] ), .B1(n3575), .B2(
        \vrf/regTable[3][104] ), .ZN(n7520) );
  AOI22D1BWP U7501 ( .A1(n3581), .A2(\vrf/regTable[0][104] ), .B1(n3594), .B2(
        \vrf/regTable[2][104] ), .ZN(n7519) );
  ND4D1BWP U7502 ( .A1(n8321), .A2(n8322), .A3(n8323), .A4(n8324), .ZN(
        scalarData1[8]) );
  AOI22D1BWP U7503 ( .A1(n8287), .A2(\srf/regTable[5][8] ), .B1(n8288), .B2(
        \srf/regTable[7][8] ), .ZN(n8324) );
  AOI22D1BWP U7504 ( .A1(n8285), .A2(\srf/regTable[4][8] ), .B1(n8286), .B2(
        \srf/regTable[6][8] ), .ZN(n8323) );
  AOI22D1BWP U7505 ( .A1(n8282), .A2(\srf/regTable[1][8] ), .B1(n8284), .B2(
        \srf/regTable[3][8] ), .ZN(n8322) );
  AOI22D1BWP U7506 ( .A1(n8278), .A2(\srf/regTable[0][8] ), .B1(n8280), .B2(
        \srf/regTable[2][8] ), .ZN(n8321) );
  AO222D1BWP U7507 ( .A1(n3669), .A2(vectorToLoad[51]), .B1(n5391), .B2(n3649), 
        .C1(n4549), .C2(n5541), .Z(N4268) );
  OAI211D1BWP U7508 ( .A1(n5335), .A2(n5509), .B(n5336), .C(n4406), .ZN(N4363)
         );
  AOI22D1BWP U7509 ( .A1(n3669), .A2(vectorToLoad[145]), .B1(n4626), .B2(n5387), .ZN(n5336) );
  AO222D1BWP U7510 ( .A1(n3640), .A2(n4548), .B1(n5526), .B2(n3667), .C1(n3669), .C2(vectorToLoad[102]), .Z(N4319) );
  NR2XD0BWP U7511 ( .A1(n4661), .A2(n5282), .ZN(n5526) );
  AO211D1BWP U7512 ( .A1(n4073), .A2(scalarData1[7]), .B(n3906), .C(n3905), 
        .Z(N4183) );
  AO22D1BWP U7513 ( .A1(n4072), .A2(vectorData1[7]), .B1(n4071), .B2(Addr[7]), 
        .Z(n3905) );
  ND4D1BWP U7514 ( .A1(n7147), .A2(n7148), .A3(n7149), .A4(n7150), .ZN(
        vectorData1[7]) );
  AOI22D1BWP U7515 ( .A1(n3576), .A2(\vrf/regTable[5][7] ), .B1(n3567), .B2(
        \vrf/regTable[7][7] ), .ZN(n7150) );
  AOI22D1BWP U7516 ( .A1(n3574), .A2(\vrf/regTable[4][7] ), .B1(n3570), .B2(
        \vrf/regTable[6][7] ), .ZN(n7149) );
  AOI22D1BWP U7517 ( .A1(n3579), .A2(\vrf/regTable[1][7] ), .B1(n3575), .B2(
        \vrf/regTable[3][7] ), .ZN(n7148) );
  AOI22D1BWP U7518 ( .A1(n3581), .A2(\vrf/regTable[0][7] ), .B1(n3572), .B2(
        \vrf/regTable[2][7] ), .ZN(n7147) );
  AOI31D1BWP U7519 ( .A1(n5069), .A2(n5068), .A3(n5070), .B(n4070), .ZN(n3906)
         );
  AOI22D1BWP U7520 ( .A1(n5231), .A2(vectorData1[119]), .B1(n5230), .B2(
        vectorData1[167]), .ZN(n5070) );
  ND4D1BWP U7521 ( .A1(n7771), .A2(n7772), .A3(n7773), .A4(n7774), .ZN(
        vectorData1[167]) );
  AOI22D1BWP U7522 ( .A1(n3576), .A2(\vrf/regTable[5][167] ), .B1(n3567), .B2(
        \vrf/regTable[7][167] ), .ZN(n7774) );
  AOI22D1BWP U7523 ( .A1(n3574), .A2(\vrf/regTable[4][167] ), .B1(n3570), .B2(
        \vrf/regTable[6][167] ), .ZN(n7773) );
  AOI22D1BWP U7524 ( .A1(n3579), .A2(\vrf/regTable[1][167] ), .B1(n3575), .B2(
        \vrf/regTable[3][167] ), .ZN(n7772) );
  AOI22D1BWP U7525 ( .A1(n3581), .A2(\vrf/regTable[0][167] ), .B1(n3572), .B2(
        \vrf/regTable[2][167] ), .ZN(n7771) );
  ND4D1BWP U7526 ( .A1(n7579), .A2(n7580), .A3(n7581), .A4(n7582), .ZN(
        vectorData1[119]) );
  AOI22D1BWP U7527 ( .A1(n3576), .A2(\vrf/regTable[5][119] ), .B1(n3567), .B2(
        \vrf/regTable[7][119] ), .ZN(n7582) );
  AOI22D1BWP U7528 ( .A1(n3574), .A2(\vrf/regTable[4][119] ), .B1(n3570), .B2(
        \vrf/regTable[6][119] ), .ZN(n7581) );
  AOI22D1BWP U7529 ( .A1(n3579), .A2(\vrf/regTable[1][119] ), .B1(n3599), .B2(
        \vrf/regTable[3][119] ), .ZN(n7580) );
  AOI22D1BWP U7530 ( .A1(n3581), .A2(\vrf/regTable[0][119] ), .B1(n3572), .B2(
        \vrf/regTable[2][119] ), .ZN(n7579) );
  AOI211XD0BWP U7531 ( .A1(n3601), .A2(vectorData1[39]), .B(n5067), .C(n5066), 
        .ZN(n5068) );
  ND4D1BWP U7532 ( .A1(n5065), .A2(n5064), .A3(n5063), .A4(n5062), .ZN(n5066)
         );
  AOI22D1BWP U7533 ( .A1(n5233), .A2(vectorData1[183]), .B1(n5184), .B2(
        vectorData1[23]), .ZN(n5062) );
  ND4D1BWP U7534 ( .A1(n7195), .A2(n7196), .A3(n7197), .A4(n7198), .ZN(
        vectorData1[23]) );
  AOI22D1BWP U7535 ( .A1(n3576), .A2(\vrf/regTable[5][23] ), .B1(n3595), .B2(
        \vrf/regTable[7][23] ), .ZN(n7198) );
  AOI22D1BWP U7536 ( .A1(n3574), .A2(\vrf/regTable[4][23] ), .B1(n3596), .B2(
        \vrf/regTable[6][23] ), .ZN(n7197) );
  AOI22D1BWP U7537 ( .A1(n3579), .A2(\vrf/regTable[1][23] ), .B1(n3599), .B2(
        \vrf/regTable[3][23] ), .ZN(n7196) );
  AOI22D1BWP U7538 ( .A1(n3581), .A2(\vrf/regTable[0][23] ), .B1(n3594), .B2(
        \vrf/regTable[2][23] ), .ZN(n7195) );
  ND4D1BWP U7539 ( .A1(n7835), .A2(n7836), .A3(n7837), .A4(n7838), .ZN(
        vectorData1[183]) );
  AOI22D1BWP U7540 ( .A1(n3576), .A2(\vrf/regTable[5][183] ), .B1(n3567), .B2(
        \vrf/regTable[7][183] ), .ZN(n7838) );
  AOI22D1BWP U7541 ( .A1(n3574), .A2(\vrf/regTable[4][183] ), .B1(n3570), .B2(
        \vrf/regTable[6][183] ), .ZN(n7837) );
  AOI22D1BWP U7542 ( .A1(n3579), .A2(\vrf/regTable[1][183] ), .B1(n3575), .B2(
        \vrf/regTable[3][183] ), .ZN(n7836) );
  AOI22D1BWP U7543 ( .A1(n3581), .A2(\vrf/regTable[0][183] ), .B1(n3572), .B2(
        \vrf/regTable[2][183] ), .ZN(n7835) );
  AOI22D1BWP U7544 ( .A1(n5226), .A2(vectorData1[135]), .B1(n5186), .B2(
        vectorData1[71]), .ZN(n5063) );
  ND4D1BWP U7545 ( .A1(n7387), .A2(n7388), .A3(n7389), .A4(n7390), .ZN(
        vectorData1[71]) );
  AOI22D1BWP U7546 ( .A1(n3576), .A2(\vrf/regTable[5][71] ), .B1(n3567), .B2(
        \vrf/regTable[7][71] ), .ZN(n7390) );
  AOI22D1BWP U7547 ( .A1(n3574), .A2(\vrf/regTable[4][71] ), .B1(n3570), .B2(
        \vrf/regTable[6][71] ), .ZN(n7389) );
  AOI22D1BWP U7548 ( .A1(n3579), .A2(\vrf/regTable[1][71] ), .B1(n3575), .B2(
        \vrf/regTable[3][71] ), .ZN(n7388) );
  AOI22D1BWP U7549 ( .A1(n3581), .A2(\vrf/regTable[0][71] ), .B1(n3572), .B2(
        \vrf/regTable[2][71] ), .ZN(n7387) );
  ND4D1BWP U7550 ( .A1(n7643), .A2(n7644), .A3(n7645), .A4(n7646), .ZN(
        vectorData1[135]) );
  AOI22D1BWP U7551 ( .A1(n3576), .A2(\vrf/regTable[5][135] ), .B1(n3567), .B2(
        \vrf/regTable[7][135] ), .ZN(n7646) );
  AOI22D1BWP U7552 ( .A1(n3574), .A2(\vrf/regTable[4][135] ), .B1(n3570), .B2(
        \vrf/regTable[6][135] ), .ZN(n7645) );
  AOI22D1BWP U7553 ( .A1(n3579), .A2(\vrf/regTable[1][135] ), .B1(n3575), .B2(
        \vrf/regTable[3][135] ), .ZN(n7644) );
  AOI22D1BWP U7554 ( .A1(n3581), .A2(\vrf/regTable[0][135] ), .B1(n3572), .B2(
        \vrf/regTable[2][135] ), .ZN(n7643) );
  AOI22D1BWP U7555 ( .A1(n5228), .A2(vectorData1[215]), .B1(n5185), .B2(
        vectorData1[87]), .ZN(n5064) );
  ND4D1BWP U7556 ( .A1(n7451), .A2(n7452), .A3(n7453), .A4(n7454), .ZN(
        vectorData1[87]) );
  AOI22D1BWP U7557 ( .A1(n7117), .A2(\vrf/regTable[5][87] ), .B1(n3567), .B2(
        \vrf/regTable[7][87] ), .ZN(n7454) );
  AOI22D1BWP U7558 ( .A1(n7115), .A2(\vrf/regTable[4][87] ), .B1(n3570), .B2(
        \vrf/regTable[6][87] ), .ZN(n7453) );
  AOI22D1BWP U7559 ( .A1(n7112), .A2(\vrf/regTable[1][87] ), .B1(n3575), .B2(
        \vrf/regTable[3][87] ), .ZN(n7452) );
  AOI22D1BWP U7560 ( .A1(n7108), .A2(\vrf/regTable[0][87] ), .B1(n3572), .B2(
        \vrf/regTable[2][87] ), .ZN(n7451) );
  ND4D1BWP U7561 ( .A1(n7963), .A2(n7964), .A3(n7965), .A4(n7966), .ZN(
        vectorData1[215]) );
  AOI22D1BWP U7562 ( .A1(n3576), .A2(\vrf/regTable[5][215] ), .B1(n3595), .B2(
        \vrf/regTable[7][215] ), .ZN(n7966) );
  AOI22D1BWP U7563 ( .A1(n3574), .A2(\vrf/regTable[4][215] ), .B1(n3596), .B2(
        \vrf/regTable[6][215] ), .ZN(n7965) );
  AOI22D1BWP U7564 ( .A1(n3579), .A2(\vrf/regTable[1][215] ), .B1(n3599), .B2(
        \vrf/regTable[3][215] ), .ZN(n7964) );
  AOI22D1BWP U7565 ( .A1(n3581), .A2(\vrf/regTable[0][215] ), .B1(n3594), .B2(
        \vrf/regTable[2][215] ), .ZN(n7963) );
  AOI22D1BWP U7566 ( .A1(n5213), .A2(vectorData1[103]), .B1(n5229), .B2(
        vectorData1[247]), .ZN(n5065) );
  ND4D1BWP U7567 ( .A1(n8091), .A2(n8092), .A3(n8093), .A4(n8094), .ZN(
        vectorData1[247]) );
  AOI22D1BWP U7568 ( .A1(n3576), .A2(\vrf/regTable[5][247] ), .B1(n7118), .B2(
        \vrf/regTable[7][247] ), .ZN(n8094) );
  AOI22D1BWP U7569 ( .A1(n3574), .A2(\vrf/regTable[4][247] ), .B1(n7116), .B2(
        \vrf/regTable[6][247] ), .ZN(n8093) );
  AOI22D1BWP U7570 ( .A1(n3579), .A2(\vrf/regTable[1][247] ), .B1(n7114), .B2(
        \vrf/regTable[3][247] ), .ZN(n8092) );
  AOI22D1BWP U7571 ( .A1(n3581), .A2(\vrf/regTable[0][247] ), .B1(n7110), .B2(
        \vrf/regTable[2][247] ), .ZN(n8091) );
  ND4D1BWP U7572 ( .A1(n7515), .A2(n7516), .A3(n7517), .A4(n7518), .ZN(
        vectorData1[103]) );
  AOI22D1BWP U7573 ( .A1(n3576), .A2(\vrf/regTable[5][103] ), .B1(n3595), .B2(
        \vrf/regTable[7][103] ), .ZN(n7518) );
  AOI22D1BWP U7574 ( .A1(n3574), .A2(\vrf/regTable[4][103] ), .B1(n3596), .B2(
        \vrf/regTable[6][103] ), .ZN(n7517) );
  AOI22D1BWP U7575 ( .A1(n3579), .A2(\vrf/regTable[1][103] ), .B1(n3575), .B2(
        \vrf/regTable[3][103] ), .ZN(n7516) );
  AOI22D1BWP U7576 ( .A1(n3581), .A2(\vrf/regTable[0][103] ), .B1(n3594), .B2(
        \vrf/regTable[2][103] ), .ZN(n7515) );
  AO22D1BWP U7577 ( .A1(n5232), .A2(vectorData1[151]), .B1(n5227), .B2(
        vectorData1[199]), .Z(n5067) );
  ND4D1BWP U7578 ( .A1(n7899), .A2(n7900), .A3(n7901), .A4(n7902), .ZN(
        vectorData1[199]) );
  AOI22D1BWP U7579 ( .A1(n3576), .A2(\vrf/regTable[5][199] ), .B1(n3567), .B2(
        \vrf/regTable[7][199] ), .ZN(n7902) );
  AOI22D1BWP U7580 ( .A1(n3574), .A2(\vrf/regTable[4][199] ), .B1(n3570), .B2(
        \vrf/regTable[6][199] ), .ZN(n7901) );
  AOI22D1BWP U7581 ( .A1(n3579), .A2(\vrf/regTable[1][199] ), .B1(n3575), .B2(
        \vrf/regTable[3][199] ), .ZN(n7900) );
  AOI22D1BWP U7582 ( .A1(n3581), .A2(\vrf/regTable[0][199] ), .B1(n3572), .B2(
        \vrf/regTable[2][199] ), .ZN(n7899) );
  ND4D1BWP U7583 ( .A1(n7707), .A2(n7708), .A3(n7709), .A4(n7710), .ZN(
        vectorData1[151]) );
  AOI22D1BWP U7584 ( .A1(n3576), .A2(\vrf/regTable[5][151] ), .B1(n3595), .B2(
        \vrf/regTable[7][151] ), .ZN(n7710) );
  AOI22D1BWP U7585 ( .A1(n3574), .A2(\vrf/regTable[4][151] ), .B1(n3596), .B2(
        \vrf/regTable[6][151] ), .ZN(n7709) );
  AOI22D1BWP U7586 ( .A1(n3579), .A2(\vrf/regTable[1][151] ), .B1(n3575), .B2(
        \vrf/regTable[3][151] ), .ZN(n7708) );
  AOI22D1BWP U7587 ( .A1(n3581), .A2(\vrf/regTable[0][151] ), .B1(n3594), .B2(
        \vrf/regTable[2][151] ), .ZN(n7707) );
  ND4D1BWP U7588 ( .A1(n7259), .A2(n7260), .A3(n7261), .A4(n7262), .ZN(
        vectorData1[39]) );
  AOI22D1BWP U7589 ( .A1(n3576), .A2(\vrf/regTable[5][39] ), .B1(n3567), .B2(
        \vrf/regTable[7][39] ), .ZN(n7262) );
  AOI22D1BWP U7590 ( .A1(n3574), .A2(\vrf/regTable[4][39] ), .B1(n3570), .B2(
        \vrf/regTable[6][39] ), .ZN(n7261) );
  AOI22D1BWP U7591 ( .A1(n3579), .A2(\vrf/regTable[1][39] ), .B1(n3575), .B2(
        \vrf/regTable[3][39] ), .ZN(n7260) );
  AOI22D1BWP U7592 ( .A1(n3581), .A2(\vrf/regTable[0][39] ), .B1(n3572), .B2(
        \vrf/regTable[2][39] ), .ZN(n7259) );
  AOI22D1BWP U7593 ( .A1(n5187), .A2(vectorData1[231]), .B1(n5188), .B2(
        vectorData1[55]), .ZN(n5069) );
  ND4D1BWP U7594 ( .A1(n7323), .A2(n7324), .A3(n7325), .A4(n7326), .ZN(
        vectorData1[55]) );
  AOI22D1BWP U7595 ( .A1(n3576), .A2(\vrf/regTable[5][55] ), .B1(n3567), .B2(
        \vrf/regTable[7][55] ), .ZN(n7326) );
  AOI22D1BWP U7596 ( .A1(n3574), .A2(\vrf/regTable[4][55] ), .B1(n3570), .B2(
        \vrf/regTable[6][55] ), .ZN(n7325) );
  AOI22D1BWP U7597 ( .A1(n3579), .A2(\vrf/regTable[1][55] ), .B1(n3575), .B2(
        \vrf/regTable[3][55] ), .ZN(n7324) );
  AOI22D1BWP U7598 ( .A1(n3581), .A2(\vrf/regTable[0][55] ), .B1(n3572), .B2(
        \vrf/regTable[2][55] ), .ZN(n7323) );
  ND4D1BWP U7599 ( .A1(n8027), .A2(n8028), .A3(n8029), .A4(n8030), .ZN(
        vectorData1[231]) );
  AOI22D1BWP U7600 ( .A1(n3576), .A2(\vrf/regTable[5][231] ), .B1(n3595), .B2(
        \vrf/regTable[7][231] ), .ZN(n8030) );
  AOI22D1BWP U7601 ( .A1(n3574), .A2(\vrf/regTable[4][231] ), .B1(n3596), .B2(
        \vrf/regTable[6][231] ), .ZN(n8029) );
  AOI22D1BWP U7602 ( .A1(n3579), .A2(\vrf/regTable[1][231] ), .B1(n3599), .B2(
        \vrf/regTable[3][231] ), .ZN(n8028) );
  AOI22D1BWP U7603 ( .A1(n3581), .A2(\vrf/regTable[0][231] ), .B1(n3594), .B2(
        \vrf/regTable[2][231] ), .ZN(n8027) );
  ND4D1BWP U7604 ( .A1(n8317), .A2(n8318), .A3(n8319), .A4(n8320), .ZN(
        scalarData1[7]) );
  AOI22D1BWP U7605 ( .A1(n8287), .A2(\srf/regTable[5][7] ), .B1(n8288), .B2(
        \srf/regTable[7][7] ), .ZN(n8320) );
  AOI22D1BWP U7606 ( .A1(n8285), .A2(\srf/regTable[4][7] ), .B1(n8286), .B2(
        \srf/regTable[6][7] ), .ZN(n8319) );
  AOI22D1BWP U7607 ( .A1(n8282), .A2(\srf/regTable[1][7] ), .B1(n8284), .B2(
        \srf/regTable[3][7] ), .ZN(n8318) );
  AOI22D1BWP U7608 ( .A1(n8278), .A2(\srf/regTable[0][7] ), .B1(n8280), .B2(
        \srf/regTable[2][7] ), .ZN(n8317) );
  OAI211D1BWP U7609 ( .A1(n5337), .A2(n5509), .B(n5338), .C(n4406), .ZN(N4364)
         );
  AOI22D1BWP U7610 ( .A1(n3669), .A2(vectorToLoad[146]), .B1(n4626), .B2(n5389), .ZN(n5338) );
  OAI211D1BWP U7611 ( .A1(n5339), .A2(n5509), .B(n5340), .C(n4406), .ZN(N4365)
         );
  AOI22D1BWP U7612 ( .A1(n3669), .A2(vectorToLoad[147]), .B1(n4626), .B2(n5391), .ZN(n5340) );
  NR2XD0BWP U7613 ( .A1(n5270), .A2(cycles[0]), .ZN(n5391) );
  AO211D1BWP U7614 ( .A1(n4073), .A2(scalarData1[6]), .B(n3857), .C(n3856), 
        .Z(N4182) );
  AO22D1BWP U7615 ( .A1(n4072), .A2(vectorData1[6]), .B1(n4071), .B2(Addr[6]), 
        .Z(n3856) );
  ND4D1BWP U7616 ( .A1(n7143), .A2(n7144), .A3(n7145), .A4(n7146), .ZN(
        vectorData1[6]) );
  AOI22D1BWP U7617 ( .A1(n3576), .A2(\vrf/regTable[5][6] ), .B1(n3567), .B2(
        \vrf/regTable[7][6] ), .ZN(n7146) );
  AOI22D1BWP U7618 ( .A1(n3574), .A2(\vrf/regTable[4][6] ), .B1(n3570), .B2(
        \vrf/regTable[6][6] ), .ZN(n7145) );
  AOI22D1BWP U7619 ( .A1(n3579), .A2(\vrf/regTable[1][6] ), .B1(n3575), .B2(
        \vrf/regTable[3][6] ), .ZN(n7144) );
  AOI22D1BWP U7620 ( .A1(n3581), .A2(\vrf/regTable[0][6] ), .B1(n3572), .B2(
        \vrf/regTable[2][6] ), .ZN(n7143) );
  AOI31D1BWP U7621 ( .A1(n5060), .A2(n5059), .A3(n5061), .B(n4070), .ZN(n3857)
         );
  AOI22D1BWP U7622 ( .A1(n5232), .A2(vectorData1[150]), .B1(n5186), .B2(
        vectorData1[70]), .ZN(n5061) );
  ND4D1BWP U7623 ( .A1(n7383), .A2(n7384), .A3(n7385), .A4(n7386), .ZN(
        vectorData1[70]) );
  AOI22D1BWP U7624 ( .A1(n3576), .A2(\vrf/regTable[5][70] ), .B1(n3595), .B2(
        \vrf/regTable[7][70] ), .ZN(n7386) );
  AOI22D1BWP U7625 ( .A1(n3574), .A2(\vrf/regTable[4][70] ), .B1(n3596), .B2(
        \vrf/regTable[6][70] ), .ZN(n7385) );
  AOI22D1BWP U7626 ( .A1(n3579), .A2(\vrf/regTable[1][70] ), .B1(n3599), .B2(
        \vrf/regTable[3][70] ), .ZN(n7384) );
  AOI22D1BWP U7627 ( .A1(n3581), .A2(\vrf/regTable[0][70] ), .B1(n3594), .B2(
        \vrf/regTable[2][70] ), .ZN(n7383) );
  ND4D1BWP U7628 ( .A1(n7703), .A2(n7704), .A3(n7705), .A4(n7706), .ZN(
        vectorData1[150]) );
  AOI22D1BWP U7629 ( .A1(n3576), .A2(\vrf/regTable[5][150] ), .B1(n3595), .B2(
        \vrf/regTable[7][150] ), .ZN(n7706) );
  AOI22D1BWP U7630 ( .A1(n3574), .A2(\vrf/regTable[4][150] ), .B1(n3596), .B2(
        \vrf/regTable[6][150] ), .ZN(n7705) );
  AOI22D1BWP U7631 ( .A1(n3579), .A2(\vrf/regTable[1][150] ), .B1(n3599), .B2(
        \vrf/regTable[3][150] ), .ZN(n7704) );
  AOI22D1BWP U7632 ( .A1(n3581), .A2(\vrf/regTable[0][150] ), .B1(n3594), .B2(
        \vrf/regTable[2][150] ), .ZN(n7703) );
  AOI211XD0BWP U7633 ( .A1(n5187), .A2(vectorData1[230]), .B(n5058), .C(n5057), 
        .ZN(n5059) );
  ND4D1BWP U7634 ( .A1(n5056), .A2(n5055), .A3(n5054), .A4(n5053), .ZN(n5057)
         );
  AOI22D1BWP U7635 ( .A1(n5229), .A2(vectorData1[246]), .B1(n5185), .B2(
        vectorData1[86]), .ZN(n5053) );
  ND4D1BWP U7636 ( .A1(n7447), .A2(n7448), .A3(n7449), .A4(n7450), .ZN(
        vectorData1[86]) );
  AOI22D1BWP U7637 ( .A1(n3576), .A2(\vrf/regTable[5][86] ), .B1(n3567), .B2(
        \vrf/regTable[7][86] ), .ZN(n7450) );
  AOI22D1BWP U7638 ( .A1(n3574), .A2(\vrf/regTable[4][86] ), .B1(n3570), .B2(
        \vrf/regTable[6][86] ), .ZN(n7449) );
  AOI22D1BWP U7639 ( .A1(n3579), .A2(\vrf/regTable[1][86] ), .B1(n3575), .B2(
        \vrf/regTable[3][86] ), .ZN(n7448) );
  AOI22D1BWP U7640 ( .A1(n3581), .A2(\vrf/regTable[0][86] ), .B1(n3572), .B2(
        \vrf/regTable[2][86] ), .ZN(n7447) );
  ND4D1BWP U7641 ( .A1(n8087), .A2(n8088), .A3(n8089), .A4(n8090), .ZN(
        vectorData1[246]) );
  AOI22D1BWP U7642 ( .A1(n3576), .A2(\vrf/regTable[5][246] ), .B1(n3595), .B2(
        \vrf/regTable[7][246] ), .ZN(n8090) );
  AOI22D1BWP U7643 ( .A1(n3574), .A2(\vrf/regTable[4][246] ), .B1(n3596), .B2(
        \vrf/regTable[6][246] ), .ZN(n8089) );
  AOI22D1BWP U7644 ( .A1(n3579), .A2(\vrf/regTable[1][246] ), .B1(n3599), .B2(
        \vrf/regTable[3][246] ), .ZN(n8088) );
  AOI22D1BWP U7645 ( .A1(n3581), .A2(\vrf/regTable[0][246] ), .B1(n3594), .B2(
        \vrf/regTable[2][246] ), .ZN(n8087) );
  AOI22D1BWP U7646 ( .A1(n3601), .A2(vectorData1[38]), .B1(n5188), .B2(
        vectorData1[54]), .ZN(n5054) );
  ND4D1BWP U7647 ( .A1(n7319), .A2(n7320), .A3(n7321), .A4(n7322), .ZN(
        vectorData1[54]) );
  AOI22D1BWP U7648 ( .A1(n3576), .A2(\vrf/regTable[5][54] ), .B1(n3567), .B2(
        \vrf/regTable[7][54] ), .ZN(n7322) );
  AOI22D1BWP U7649 ( .A1(n3574), .A2(\vrf/regTable[4][54] ), .B1(n3570), .B2(
        \vrf/regTable[6][54] ), .ZN(n7321) );
  AOI22D1BWP U7650 ( .A1(n3579), .A2(\vrf/regTable[1][54] ), .B1(n3575), .B2(
        \vrf/regTable[3][54] ), .ZN(n7320) );
  AOI22D1BWP U7651 ( .A1(n3581), .A2(\vrf/regTable[0][54] ), .B1(n3572), .B2(
        \vrf/regTable[2][54] ), .ZN(n7319) );
  ND4D1BWP U7652 ( .A1(n7255), .A2(n7256), .A3(n7257), .A4(n7258), .ZN(
        vectorData1[38]) );
  AOI22D1BWP U7653 ( .A1(n3576), .A2(\vrf/regTable[5][38] ), .B1(n3595), .B2(
        \vrf/regTable[7][38] ), .ZN(n7258) );
  AOI22D1BWP U7654 ( .A1(n3574), .A2(\vrf/regTable[4][38] ), .B1(n3596), .B2(
        \vrf/regTable[6][38] ), .ZN(n7257) );
  AOI22D1BWP U7655 ( .A1(n3579), .A2(\vrf/regTable[1][38] ), .B1(n3599), .B2(
        \vrf/regTable[3][38] ), .ZN(n7256) );
  AOI22D1BWP U7656 ( .A1(n3581), .A2(\vrf/regTable[0][38] ), .B1(n3594), .B2(
        \vrf/regTable[2][38] ), .ZN(n7255) );
  AOI22D1BWP U7657 ( .A1(n5213), .A2(vectorData1[102]), .B1(n5228), .B2(
        vectorData1[214]), .ZN(n5055) );
  ND4D1BWP U7658 ( .A1(n7959), .A2(n7960), .A3(n7961), .A4(n7962), .ZN(
        vectorData1[214]) );
  AOI22D1BWP U7659 ( .A1(n3576), .A2(\vrf/regTable[5][214] ), .B1(n3595), .B2(
        \vrf/regTable[7][214] ), .ZN(n7962) );
  AOI22D1BWP U7660 ( .A1(n3574), .A2(\vrf/regTable[4][214] ), .B1(n3596), .B2(
        \vrf/regTable[6][214] ), .ZN(n7961) );
  AOI22D1BWP U7661 ( .A1(n3579), .A2(\vrf/regTable[1][214] ), .B1(n3599), .B2(
        \vrf/regTable[3][214] ), .ZN(n7960) );
  AOI22D1BWP U7662 ( .A1(n3581), .A2(\vrf/regTable[0][214] ), .B1(n3594), .B2(
        \vrf/regTable[2][214] ), .ZN(n7959) );
  ND4D1BWP U7663 ( .A1(n7511), .A2(n7512), .A3(n7513), .A4(n7514), .ZN(
        vectorData1[102]) );
  AOI22D1BWP U7664 ( .A1(n3576), .A2(\vrf/regTable[5][102] ), .B1(n3595), .B2(
        \vrf/regTable[7][102] ), .ZN(n7514) );
  AOI22D1BWP U7665 ( .A1(n3574), .A2(\vrf/regTable[4][102] ), .B1(n3596), .B2(
        \vrf/regTable[6][102] ), .ZN(n7513) );
  AOI22D1BWP U7666 ( .A1(n3579), .A2(\vrf/regTable[1][102] ), .B1(n3575), .B2(
        \vrf/regTable[3][102] ), .ZN(n7512) );
  AOI22D1BWP U7667 ( .A1(n3581), .A2(\vrf/regTable[0][102] ), .B1(n3594), .B2(
        \vrf/regTable[2][102] ), .ZN(n7511) );
  AOI22D1BWP U7668 ( .A1(n5226), .A2(vectorData1[134]), .B1(n5231), .B2(
        vectorData1[118]), .ZN(n5056) );
  ND4D1BWP U7669 ( .A1(n7575), .A2(n7576), .A3(n7577), .A4(n7578), .ZN(
        vectorData1[118]) );
  AOI22D1BWP U7670 ( .A1(n3576), .A2(\vrf/regTable[5][118] ), .B1(n3595), .B2(
        \vrf/regTable[7][118] ), .ZN(n7578) );
  AOI22D1BWP U7671 ( .A1(n3574), .A2(\vrf/regTable[4][118] ), .B1(n3596), .B2(
        \vrf/regTable[6][118] ), .ZN(n7577) );
  AOI22D1BWP U7672 ( .A1(n3579), .A2(\vrf/regTable[1][118] ), .B1(n3575), .B2(
        \vrf/regTable[3][118] ), .ZN(n7576) );
  AOI22D1BWP U7673 ( .A1(n3581), .A2(\vrf/regTable[0][118] ), .B1(n3594), .B2(
        \vrf/regTable[2][118] ), .ZN(n7575) );
  ND4D1BWP U7674 ( .A1(n7639), .A2(n7640), .A3(n7641), .A4(n7642), .ZN(
        vectorData1[134]) );
  AOI22D1BWP U7675 ( .A1(n3576), .A2(\vrf/regTable[5][134] ), .B1(n3567), .B2(
        \vrf/regTable[7][134] ), .ZN(n7642) );
  AOI22D1BWP U7676 ( .A1(n3574), .A2(\vrf/regTable[4][134] ), .B1(n3570), .B2(
        \vrf/regTable[6][134] ), .ZN(n7641) );
  AOI22D1BWP U7677 ( .A1(n3579), .A2(\vrf/regTable[1][134] ), .B1(n3599), .B2(
        \vrf/regTable[3][134] ), .ZN(n7640) );
  AOI22D1BWP U7678 ( .A1(n3581), .A2(\vrf/regTable[0][134] ), .B1(n3572), .B2(
        \vrf/regTable[2][134] ), .ZN(n7639) );
  AO22D1BWP U7679 ( .A1(n5230), .A2(vectorData1[166]), .B1(n5227), .B2(
        vectorData1[198]), .Z(n5058) );
  ND4D1BWP U7680 ( .A1(n7895), .A2(n7896), .A3(n7897), .A4(n7898), .ZN(
        vectorData1[198]) );
  AOI22D1BWP U7681 ( .A1(n3576), .A2(\vrf/regTable[5][198] ), .B1(n3595), .B2(
        \vrf/regTable[7][198] ), .ZN(n7898) );
  AOI22D1BWP U7682 ( .A1(n3574), .A2(\vrf/regTable[4][198] ), .B1(n3596), .B2(
        \vrf/regTable[6][198] ), .ZN(n7897) );
  AOI22D1BWP U7683 ( .A1(n3579), .A2(\vrf/regTable[1][198] ), .B1(n3599), .B2(
        \vrf/regTable[3][198] ), .ZN(n7896) );
  AOI22D1BWP U7684 ( .A1(n3581), .A2(\vrf/regTable[0][198] ), .B1(n3594), .B2(
        \vrf/regTable[2][198] ), .ZN(n7895) );
  ND4D1BWP U7685 ( .A1(n7767), .A2(n7768), .A3(n7769), .A4(n7770), .ZN(
        vectorData1[166]) );
  AOI22D1BWP U7686 ( .A1(n3576), .A2(\vrf/regTable[5][166] ), .B1(n3567), .B2(
        \vrf/regTable[7][166] ), .ZN(n7770) );
  AOI22D1BWP U7687 ( .A1(n3574), .A2(\vrf/regTable[4][166] ), .B1(n3570), .B2(
        \vrf/regTable[6][166] ), .ZN(n7769) );
  AOI22D1BWP U7688 ( .A1(n3579), .A2(\vrf/regTable[1][166] ), .B1(n3575), .B2(
        \vrf/regTable[3][166] ), .ZN(n7768) );
  AOI22D1BWP U7689 ( .A1(n3581), .A2(\vrf/regTable[0][166] ), .B1(n3572), .B2(
        \vrf/regTable[2][166] ), .ZN(n7767) );
  ND4D1BWP U7690 ( .A1(n8023), .A2(n8024), .A3(n8025), .A4(n8026), .ZN(
        vectorData1[230]) );
  AOI22D1BWP U7691 ( .A1(n3576), .A2(\vrf/regTable[5][230] ), .B1(n3567), .B2(
        \vrf/regTable[7][230] ), .ZN(n8026) );
  AOI22D1BWP U7692 ( .A1(n3574), .A2(\vrf/regTable[4][230] ), .B1(n3570), .B2(
        \vrf/regTable[6][230] ), .ZN(n8025) );
  AOI22D1BWP U7693 ( .A1(n3579), .A2(\vrf/regTable[1][230] ), .B1(n3575), .B2(
        \vrf/regTable[3][230] ), .ZN(n8024) );
  AOI22D1BWP U7694 ( .A1(n3581), .A2(\vrf/regTable[0][230] ), .B1(n3572), .B2(
        \vrf/regTable[2][230] ), .ZN(n8023) );
  AOI22D1BWP U7695 ( .A1(n5233), .A2(vectorData1[182]), .B1(n5184), .B2(
        vectorData1[22]), .ZN(n5060) );
  ND4D1BWP U7696 ( .A1(n7191), .A2(n7192), .A3(n7193), .A4(n7194), .ZN(
        vectorData1[22]) );
  AOI22D1BWP U7697 ( .A1(n3576), .A2(\vrf/regTable[5][22] ), .B1(n3567), .B2(
        \vrf/regTable[7][22] ), .ZN(n7194) );
  AOI22D1BWP U7698 ( .A1(n3574), .A2(\vrf/regTable[4][22] ), .B1(n3570), .B2(
        \vrf/regTable[6][22] ), .ZN(n7193) );
  AOI22D1BWP U7699 ( .A1(n3579), .A2(\vrf/regTable[1][22] ), .B1(n3575), .B2(
        \vrf/regTable[3][22] ), .ZN(n7192) );
  AOI22D1BWP U7700 ( .A1(n3581), .A2(\vrf/regTable[0][22] ), .B1(n3572), .B2(
        \vrf/regTable[2][22] ), .ZN(n7191) );
  ND4D1BWP U7701 ( .A1(n7831), .A2(n7832), .A3(n7833), .A4(n7834), .ZN(
        vectorData1[182]) );
  AOI22D1BWP U7702 ( .A1(n3576), .A2(\vrf/regTable[5][182] ), .B1(n3567), .B2(
        \vrf/regTable[7][182] ), .ZN(n7834) );
  AOI22D1BWP U7703 ( .A1(n3574), .A2(\vrf/regTable[4][182] ), .B1(n3570), .B2(
        \vrf/regTable[6][182] ), .ZN(n7833) );
  AOI22D1BWP U7704 ( .A1(n3579), .A2(\vrf/regTable[1][182] ), .B1(n3575), .B2(
        \vrf/regTable[3][182] ), .ZN(n7832) );
  AOI22D1BWP U7705 ( .A1(n3581), .A2(\vrf/regTable[0][182] ), .B1(n3572), .B2(
        \vrf/regTable[2][182] ), .ZN(n7831) );
  ND4D1BWP U7706 ( .A1(n8313), .A2(n8314), .A3(n8315), .A4(n8316), .ZN(
        scalarData1[6]) );
  AOI22D1BWP U7707 ( .A1(n8287), .A2(\srf/regTable[5][6] ), .B1(n8288), .B2(
        \srf/regTable[7][6] ), .ZN(n8316) );
  AOI22D1BWP U7708 ( .A1(n8285), .A2(\srf/regTable[4][6] ), .B1(n8286), .B2(
        \srf/regTable[6][6] ), .ZN(n8315) );
  AOI22D1BWP U7709 ( .A1(n8282), .A2(\srf/regTable[1][6] ), .B1(n8284), .B2(
        \srf/regTable[3][6] ), .ZN(n8314) );
  AOI22D1BWP U7710 ( .A1(n8278), .A2(\srf/regTable[0][6] ), .B1(n8280), .B2(
        \srf/regTable[2][6] ), .ZN(n8313) );
  OAI211D1BWP U7711 ( .A1(n5476), .A2(n4405), .B(n5343), .C(n4535), .ZN(N4366)
         );
  AOI22D1BWP U7712 ( .A1(n3669), .A2(vectorToLoad[148]), .B1(n4627), .B2(n5342), .ZN(n5343) );
  NR2XD0BWP U7713 ( .A1(n5334), .A2(n4665), .ZN(n5342) );
  NR2XD0BWP U7714 ( .A1(n5271), .A2(cycles[0]), .ZN(n5341) );
  AO222D1BWP U7715 ( .A1(n3668), .A2(vectorToLoad[50]), .B1(n5389), .B2(n3649), 
        .C1(n4549), .C2(n5540), .Z(N4267) );
  NR2XD0BWP U7716 ( .A1(n5269), .A2(cycles[0]), .ZN(n5389) );
  OAI211D1BWP U7717 ( .A1(n5344), .A2(n5509), .B(n5345), .C(n4406), .ZN(N4367)
         );
  AOI22D1BWP U7718 ( .A1(n3669), .A2(vectorToLoad[149]), .B1(n4626), .B2(n5394), .ZN(n5345) );
  NR2XD0BWP U7719 ( .A1(n5272), .A2(cycles[0]), .ZN(n5394) );
  AO211D1BWP U7720 ( .A1(n4073), .A2(scalarData1[5]), .B(n3847), .C(n3846), 
        .Z(N4181) );
  AO22D1BWP U7721 ( .A1(n4072), .A2(vectorData1[5]), .B1(n4071), .B2(Addr[5]), 
        .Z(n3846) );
  ND4D1BWP U7722 ( .A1(n7139), .A2(n7140), .A3(n7141), .A4(n7142), .ZN(
        vectorData1[5]) );
  AOI22D1BWP U7723 ( .A1(n3576), .A2(\vrf/regTable[5][5] ), .B1(n3567), .B2(
        \vrf/regTable[7][5] ), .ZN(n7142) );
  AOI22D1BWP U7724 ( .A1(n3574), .A2(\vrf/regTable[4][5] ), .B1(n3570), .B2(
        \vrf/regTable[6][5] ), .ZN(n7141) );
  AOI22D1BWP U7725 ( .A1(n3579), .A2(\vrf/regTable[1][5] ), .B1(n3575), .B2(
        \vrf/regTable[3][5] ), .ZN(n7140) );
  AOI22D1BWP U7726 ( .A1(n3581), .A2(\vrf/regTable[0][5] ), .B1(n3572), .B2(
        \vrf/regTable[2][5] ), .ZN(n7139) );
  AOI31D1BWP U7727 ( .A1(n5051), .A2(n5050), .A3(n5052), .B(n4070), .ZN(n3847)
         );
  AOI22D1BWP U7728 ( .A1(n3601), .A2(vectorData1[37]), .B1(n5230), .B2(
        vectorData1[165]), .ZN(n5052) );
  ND4D1BWP U7729 ( .A1(n7763), .A2(n7764), .A3(n7765), .A4(n7766), .ZN(
        vectorData1[165]) );
  AOI22D1BWP U7730 ( .A1(n3576), .A2(\vrf/regTable[5][165] ), .B1(n3567), .B2(
        \vrf/regTable[7][165] ), .ZN(n7766) );
  AOI22D1BWP U7731 ( .A1(n3574), .A2(\vrf/regTable[4][165] ), .B1(n3570), .B2(
        \vrf/regTable[6][165] ), .ZN(n7765) );
  AOI22D1BWP U7732 ( .A1(n3579), .A2(\vrf/regTable[1][165] ), .B1(n3575), .B2(
        \vrf/regTable[3][165] ), .ZN(n7764) );
  AOI22D1BWP U7733 ( .A1(n3581), .A2(\vrf/regTable[0][165] ), .B1(n3572), .B2(
        \vrf/regTable[2][165] ), .ZN(n7763) );
  ND4D1BWP U7734 ( .A1(n7251), .A2(n7252), .A3(n7253), .A4(n7254), .ZN(
        vectorData1[37]) );
  AOI22D1BWP U7735 ( .A1(n3576), .A2(\vrf/regTable[5][37] ), .B1(n3595), .B2(
        \vrf/regTable[7][37] ), .ZN(n7254) );
  AOI22D1BWP U7736 ( .A1(n3574), .A2(\vrf/regTable[4][37] ), .B1(n3596), .B2(
        \vrf/regTable[6][37] ), .ZN(n7253) );
  AOI22D1BWP U7737 ( .A1(n3579), .A2(\vrf/regTable[1][37] ), .B1(n3599), .B2(
        \vrf/regTable[3][37] ), .ZN(n7252) );
  AOI22D1BWP U7738 ( .A1(n3581), .A2(\vrf/regTable[0][37] ), .B1(n3594), .B2(
        \vrf/regTable[2][37] ), .ZN(n7251) );
  AOI211XD0BWP U7739 ( .A1(n5226), .A2(vectorData1[133]), .B(n5049), .C(n5048), 
        .ZN(n5050) );
  ND4D1BWP U7740 ( .A1(n5047), .A2(n5046), .A3(n5045), .A4(n5044), .ZN(n5048)
         );
  AOI22D1BWP U7741 ( .A1(n5185), .A2(vectorData1[85]), .B1(n5188), .B2(
        vectorData1[53]), .ZN(n5044) );
  ND4D1BWP U7742 ( .A1(n7315), .A2(n7316), .A3(n7317), .A4(n7318), .ZN(
        vectorData1[53]) );
  AOI22D1BWP U7743 ( .A1(n3576), .A2(\vrf/regTable[5][53] ), .B1(n3567), .B2(
        \vrf/regTable[7][53] ), .ZN(n7318) );
  AOI22D1BWP U7744 ( .A1(n3574), .A2(\vrf/regTable[4][53] ), .B1(n3570), .B2(
        \vrf/regTable[6][53] ), .ZN(n7317) );
  AOI22D1BWP U7745 ( .A1(n3579), .A2(\vrf/regTable[1][53] ), .B1(n3575), .B2(
        \vrf/regTable[3][53] ), .ZN(n7316) );
  AOI22D1BWP U7746 ( .A1(n3581), .A2(\vrf/regTable[0][53] ), .B1(n3572), .B2(
        \vrf/regTable[2][53] ), .ZN(n7315) );
  ND4D1BWP U7747 ( .A1(n7443), .A2(n7444), .A3(n7445), .A4(n7446), .ZN(
        vectorData1[85]) );
  AOI22D1BWP U7748 ( .A1(n3576), .A2(\vrf/regTable[5][85] ), .B1(n3567), .B2(
        \vrf/regTable[7][85] ), .ZN(n7446) );
  AOI22D1BWP U7749 ( .A1(n3574), .A2(\vrf/regTable[4][85] ), .B1(n3570), .B2(
        \vrf/regTable[6][85] ), .ZN(n7445) );
  AOI22D1BWP U7750 ( .A1(n3579), .A2(\vrf/regTable[1][85] ), .B1(n3575), .B2(
        \vrf/regTable[3][85] ), .ZN(n7444) );
  AOI22D1BWP U7751 ( .A1(n3581), .A2(\vrf/regTable[0][85] ), .B1(n3572), .B2(
        \vrf/regTable[2][85] ), .ZN(n7443) );
  AOI22D1BWP U7752 ( .A1(n5213), .A2(vectorData1[101]), .B1(n5228), .B2(
        vectorData1[213]), .ZN(n5045) );
  ND4D1BWP U7753 ( .A1(n7955), .A2(n7956), .A3(n7957), .A4(n7958), .ZN(
        vectorData1[213]) );
  AOI22D1BWP U7754 ( .A1(n3576), .A2(\vrf/regTable[5][213] ), .B1(n3595), .B2(
        \vrf/regTable[7][213] ), .ZN(n7958) );
  AOI22D1BWP U7755 ( .A1(n3574), .A2(\vrf/regTable[4][213] ), .B1(n3596), .B2(
        \vrf/regTable[6][213] ), .ZN(n7957) );
  AOI22D1BWP U7756 ( .A1(n3579), .A2(\vrf/regTable[1][213] ), .B1(n3599), .B2(
        \vrf/regTable[3][213] ), .ZN(n7956) );
  AOI22D1BWP U7757 ( .A1(n3581), .A2(\vrf/regTable[0][213] ), .B1(n3594), .B2(
        \vrf/regTable[2][213] ), .ZN(n7955) );
  ND4D1BWP U7758 ( .A1(n7507), .A2(n7508), .A3(n7509), .A4(n7510), .ZN(
        vectorData1[101]) );
  AOI22D1BWP U7759 ( .A1(n7117), .A2(\vrf/regTable[5][101] ), .B1(n3595), .B2(
        \vrf/regTable[7][101] ), .ZN(n7510) );
  AOI22D1BWP U7760 ( .A1(n7115), .A2(\vrf/regTable[4][101] ), .B1(n3596), .B2(
        \vrf/regTable[6][101] ), .ZN(n7509) );
  AOI22D1BWP U7761 ( .A1(n7112), .A2(\vrf/regTable[1][101] ), .B1(n3599), .B2(
        \vrf/regTable[3][101] ), .ZN(n7508) );
  AOI22D1BWP U7762 ( .A1(n7108), .A2(\vrf/regTable[0][101] ), .B1(n3594), .B2(
        \vrf/regTable[2][101] ), .ZN(n7507) );
  AOI22D1BWP U7763 ( .A1(n5232), .A2(vectorData1[149]), .B1(n5227), .B2(
        vectorData1[197]), .ZN(n5046) );
  ND4D1BWP U7764 ( .A1(n7891), .A2(n7892), .A3(n7893), .A4(n7894), .ZN(
        vectorData1[197]) );
  AOI22D1BWP U7765 ( .A1(n3576), .A2(\vrf/regTable[5][197] ), .B1(n7118), .B2(
        \vrf/regTable[7][197] ), .ZN(n7894) );
  AOI22D1BWP U7766 ( .A1(n3574), .A2(\vrf/regTable[4][197] ), .B1(n7116), .B2(
        \vrf/regTable[6][197] ), .ZN(n7893) );
  AOI22D1BWP U7767 ( .A1(n3579), .A2(\vrf/regTable[1][197] ), .B1(n7114), .B2(
        \vrf/regTable[3][197] ), .ZN(n7892) );
  AOI22D1BWP U7768 ( .A1(n3581), .A2(\vrf/regTable[0][197] ), .B1(n7110), .B2(
        \vrf/regTable[2][197] ), .ZN(n7891) );
  ND4D1BWP U7769 ( .A1(n7699), .A2(n7700), .A3(n7701), .A4(n7702), .ZN(
        vectorData1[149]) );
  AOI22D1BWP U7770 ( .A1(n3576), .A2(\vrf/regTable[5][149] ), .B1(n3595), .B2(
        \vrf/regTable[7][149] ), .ZN(n7702) );
  AOI22D1BWP U7771 ( .A1(n3574), .A2(\vrf/regTable[4][149] ), .B1(n3596), .B2(
        \vrf/regTable[6][149] ), .ZN(n7701) );
  AOI22D1BWP U7772 ( .A1(n3579), .A2(\vrf/regTable[1][149] ), .B1(n3575), .B2(
        \vrf/regTable[3][149] ), .ZN(n7700) );
  AOI22D1BWP U7773 ( .A1(n3581), .A2(\vrf/regTable[0][149] ), .B1(n3594), .B2(
        \vrf/regTable[2][149] ), .ZN(n7699) );
  AOI22D1BWP U7774 ( .A1(n5229), .A2(vectorData1[245]), .B1(n5184), .B2(
        vectorData1[21]), .ZN(n5047) );
  ND4D1BWP U7775 ( .A1(n7187), .A2(n7188), .A3(n7189), .A4(n7190), .ZN(
        vectorData1[21]) );
  AOI22D1BWP U7776 ( .A1(n3576), .A2(\vrf/regTable[5][21] ), .B1(n3595), .B2(
        \vrf/regTable[7][21] ), .ZN(n7190) );
  AOI22D1BWP U7777 ( .A1(n3574), .A2(\vrf/regTable[4][21] ), .B1(n3596), .B2(
        \vrf/regTable[6][21] ), .ZN(n7189) );
  AOI22D1BWP U7778 ( .A1(n3579), .A2(\vrf/regTable[1][21] ), .B1(n3599), .B2(
        \vrf/regTable[3][21] ), .ZN(n7188) );
  AOI22D1BWP U7779 ( .A1(n3581), .A2(\vrf/regTable[0][21] ), .B1(n3594), .B2(
        \vrf/regTable[2][21] ), .ZN(n7187) );
  ND4D1BWP U7780 ( .A1(n8083), .A2(n8084), .A3(n8085), .A4(n8086), .ZN(
        vectorData1[245]) );
  AOI22D1BWP U7781 ( .A1(n3576), .A2(\vrf/regTable[5][245] ), .B1(n3595), .B2(
        \vrf/regTable[7][245] ), .ZN(n8086) );
  AOI22D1BWP U7782 ( .A1(n3574), .A2(\vrf/regTable[4][245] ), .B1(n3596), .B2(
        \vrf/regTable[6][245] ), .ZN(n8085) );
  AOI22D1BWP U7783 ( .A1(n3579), .A2(\vrf/regTable[1][245] ), .B1(n3599), .B2(
        \vrf/regTable[3][245] ), .ZN(n8084) );
  AOI22D1BWP U7784 ( .A1(n3581), .A2(\vrf/regTable[0][245] ), .B1(n3594), .B2(
        \vrf/regTable[2][245] ), .ZN(n8083) );
  AO22D1BWP U7785 ( .A1(n5187), .A2(vectorData1[229]), .B1(n5186), .B2(
        vectorData1[69]), .Z(n5049) );
  ND4D1BWP U7786 ( .A1(n7379), .A2(n7380), .A3(n7381), .A4(n7382), .ZN(
        vectorData1[69]) );
  AOI22D1BWP U7787 ( .A1(n3576), .A2(\vrf/regTable[5][69] ), .B1(n3595), .B2(
        \vrf/regTable[7][69] ), .ZN(n7382) );
  AOI22D1BWP U7788 ( .A1(n3574), .A2(\vrf/regTable[4][69] ), .B1(n3596), .B2(
        \vrf/regTable[6][69] ), .ZN(n7381) );
  AOI22D1BWP U7789 ( .A1(n3579), .A2(\vrf/regTable[1][69] ), .B1(n3599), .B2(
        \vrf/regTable[3][69] ), .ZN(n7380) );
  AOI22D1BWP U7790 ( .A1(n3581), .A2(\vrf/regTable[0][69] ), .B1(n3594), .B2(
        \vrf/regTable[2][69] ), .ZN(n7379) );
  ND4D1BWP U7791 ( .A1(n8019), .A2(n8020), .A3(n8021), .A4(n8022), .ZN(
        vectorData1[229]) );
  AOI22D1BWP U7792 ( .A1(n3576), .A2(\vrf/regTable[5][229] ), .B1(n3567), .B2(
        \vrf/regTable[7][229] ), .ZN(n8022) );
  AOI22D1BWP U7793 ( .A1(n3574), .A2(\vrf/regTable[4][229] ), .B1(n3570), .B2(
        \vrf/regTable[6][229] ), .ZN(n8021) );
  AOI22D1BWP U7794 ( .A1(n3579), .A2(\vrf/regTable[1][229] ), .B1(n3575), .B2(
        \vrf/regTable[3][229] ), .ZN(n8020) );
  AOI22D1BWP U7795 ( .A1(n3581), .A2(\vrf/regTable[0][229] ), .B1(n3572), .B2(
        \vrf/regTable[2][229] ), .ZN(n8019) );
  ND4D1BWP U7796 ( .A1(n7635), .A2(n7636), .A3(n7637), .A4(n7638), .ZN(
        vectorData1[133]) );
  AOI22D1BWP U7797 ( .A1(n3576), .A2(\vrf/regTable[5][133] ), .B1(n3567), .B2(
        \vrf/regTable[7][133] ), .ZN(n7638) );
  AOI22D1BWP U7798 ( .A1(n3574), .A2(\vrf/regTable[4][133] ), .B1(n3570), .B2(
        \vrf/regTable[6][133] ), .ZN(n7637) );
  AOI22D1BWP U7799 ( .A1(n3579), .A2(\vrf/regTable[1][133] ), .B1(n3575), .B2(
        \vrf/regTable[3][133] ), .ZN(n7636) );
  AOI22D1BWP U7800 ( .A1(n3581), .A2(\vrf/regTable[0][133] ), .B1(n3572), .B2(
        \vrf/regTable[2][133] ), .ZN(n7635) );
  AOI22D1BWP U7801 ( .A1(n5231), .A2(vectorData1[117]), .B1(n5233), .B2(
        vectorData1[181]), .ZN(n5051) );
  ND4D1BWP U7802 ( .A1(n7827), .A2(n7828), .A3(n7829), .A4(n7830), .ZN(
        vectorData1[181]) );
  AOI22D1BWP U7803 ( .A1(n3576), .A2(\vrf/regTable[5][181] ), .B1(n3595), .B2(
        \vrf/regTable[7][181] ), .ZN(n7830) );
  AOI22D1BWP U7804 ( .A1(n3574), .A2(\vrf/regTable[4][181] ), .B1(n3596), .B2(
        \vrf/regTable[6][181] ), .ZN(n7829) );
  AOI22D1BWP U7805 ( .A1(n3579), .A2(\vrf/regTable[1][181] ), .B1(n3599), .B2(
        \vrf/regTable[3][181] ), .ZN(n7828) );
  AOI22D1BWP U7806 ( .A1(n3581), .A2(\vrf/regTable[0][181] ), .B1(n3594), .B2(
        \vrf/regTable[2][181] ), .ZN(n7827) );
  ND4D1BWP U7807 ( .A1(n7571), .A2(n7572), .A3(n7573), .A4(n7574), .ZN(
        vectorData1[117]) );
  AOI22D1BWP U7808 ( .A1(n3576), .A2(\vrf/regTable[5][117] ), .B1(n3567), .B2(
        \vrf/regTable[7][117] ), .ZN(n7574) );
  AOI22D1BWP U7809 ( .A1(n3574), .A2(\vrf/regTable[4][117] ), .B1(n3570), .B2(
        \vrf/regTable[6][117] ), .ZN(n7573) );
  AOI22D1BWP U7810 ( .A1(n3579), .A2(\vrf/regTable[1][117] ), .B1(n3599), .B2(
        \vrf/regTable[3][117] ), .ZN(n7572) );
  AOI22D1BWP U7811 ( .A1(n3581), .A2(\vrf/regTable[0][117] ), .B1(n3572), .B2(
        \vrf/regTable[2][117] ), .ZN(n7571) );
  ND4D1BWP U7812 ( .A1(n8309), .A2(n8310), .A3(n8311), .A4(n8312), .ZN(
        scalarData1[5]) );
  AOI22D1BWP U7813 ( .A1(n8287), .A2(\srf/regTable[5][5] ), .B1(n8288), .B2(
        \srf/regTable[7][5] ), .ZN(n8312) );
  AOI22D1BWP U7814 ( .A1(n8285), .A2(\srf/regTable[4][5] ), .B1(n8286), .B2(
        \srf/regTable[6][5] ), .ZN(n8311) );
  AOI22D1BWP U7815 ( .A1(n8282), .A2(\srf/regTable[1][5] ), .B1(n8284), .B2(
        \srf/regTable[3][5] ), .ZN(n8310) );
  AOI22D1BWP U7816 ( .A1(n8278), .A2(\srf/regTable[0][5] ), .B1(n8280), .B2(
        \srf/regTable[2][5] ), .ZN(n8309) );
  OAI211D1BWP U7817 ( .A1(n5346), .A2(n5509), .B(n5347), .C(n4406), .ZN(N4368)
         );
  AOI22D1BWP U7818 ( .A1(n3669), .A2(vectorToLoad[150]), .B1(n4626), .B2(n5396), .ZN(n5347) );
  NR2XD0BWP U7819 ( .A1(n5273), .A2(cycles[0]), .ZN(n5396) );
  AO222D1BWP U7820 ( .A1(n3668), .A2(vectorToLoad[49]), .B1(n4549), .B2(n5539), 
        .C1(n3649), .C2(n5387), .Z(N4266) );
  NR2XD0BWP U7821 ( .A1(n5268), .A2(cycles[0]), .ZN(n5387) );
  OAI211D1BWP U7822 ( .A1(n5348), .A2(n5509), .B(n5349), .C(n4406), .ZN(N4369)
         );
  AOI22D1BWP U7823 ( .A1(n3669), .A2(vectorToLoad[151]), .B1(n4626), .B2(n5398), .ZN(n5349) );
  NR2XD0BWP U7824 ( .A1(n5274), .A2(cycles[0]), .ZN(n5398) );
  OAI211D1BWP U7825 ( .A1(n3833), .A2(n4070), .B(n3832), .C(n3831), .ZN(N4180)
         );
  ND4D1BWP U7826 ( .A1(n8305), .A2(n8306), .A3(n8307), .A4(n8308), .ZN(
        scalarData1[4]) );
  AOI22D1BWP U7827 ( .A1(n8287), .A2(\srf/regTable[5][4] ), .B1(n8288), .B2(
        \srf/regTable[7][4] ), .ZN(n8308) );
  AOI22D1BWP U7828 ( .A1(n8285), .A2(\srf/regTable[4][4] ), .B1(n8286), .B2(
        \srf/regTable[6][4] ), .ZN(n8307) );
  AOI22D1BWP U7829 ( .A1(n8282), .A2(\srf/regTable[1][4] ), .B1(n8284), .B2(
        \srf/regTable[3][4] ), .ZN(n8306) );
  AOI22D1BWP U7830 ( .A1(n8278), .A2(\srf/regTable[0][4] ), .B1(n8280), .B2(
        \srf/regTable[2][4] ), .ZN(n8305) );
  AOI22D1BWP U7831 ( .A1(n4072), .A2(vectorData1[4]), .B1(n4071), .B2(Addr[4]), 
        .ZN(n3832) );
  ND4D1BWP U7832 ( .A1(n7135), .A2(n7136), .A3(n7137), .A4(n7138), .ZN(
        vectorData1[4]) );
  AOI22D1BWP U7833 ( .A1(n3576), .A2(\vrf/regTable[5][4] ), .B1(n3595), .B2(
        \vrf/regTable[7][4] ), .ZN(n7138) );
  AOI22D1BWP U7834 ( .A1(n3574), .A2(\vrf/regTable[4][4] ), .B1(n3596), .B2(
        \vrf/regTable[6][4] ), .ZN(n7137) );
  AOI22D1BWP U7835 ( .A1(n3579), .A2(\vrf/regTable[1][4] ), .B1(n3599), .B2(
        \vrf/regTable[3][4] ), .ZN(n7136) );
  AOI22D1BWP U7836 ( .A1(n3581), .A2(\vrf/regTable[0][4] ), .B1(n3594), .B2(
        \vrf/regTable[2][4] ), .ZN(n7135) );
  AOI211XD0BWP U7837 ( .A1(n5187), .A2(vectorData1[228]), .B(n3829), .C(n3828), 
        .ZN(n3833) );
  IND3D1BWP U7838 ( .A1(n5040), .B1(n5042), .B2(n3827), .ZN(n3828) );
  ND4D1BWP U7839 ( .A1(n7375), .A2(n7376), .A3(n7377), .A4(n7378), .ZN(
        vectorData1[68]) );
  AOI22D1BWP U7840 ( .A1(n3576), .A2(\vrf/regTable[5][68] ), .B1(n3567), .B2(
        \vrf/regTable[7][68] ), .ZN(n7378) );
  AOI22D1BWP U7841 ( .A1(n3574), .A2(\vrf/regTable[4][68] ), .B1(n3570), .B2(
        \vrf/regTable[6][68] ), .ZN(n7377) );
  AOI22D1BWP U7842 ( .A1(n3579), .A2(\vrf/regTable[1][68] ), .B1(n3575), .B2(
        \vrf/regTable[3][68] ), .ZN(n7376) );
  AOI22D1BWP U7843 ( .A1(n3581), .A2(\vrf/regTable[0][68] ), .B1(n3572), .B2(
        \vrf/regTable[2][68] ), .ZN(n7375) );
  AOI22D1BWP U7844 ( .A1(n5228), .A2(vectorData1[212]), .B1(n5188), .B2(
        vectorData1[52]), .ZN(n5042) );
  ND4D1BWP U7845 ( .A1(n7311), .A2(n7312), .A3(n7313), .A4(n7314), .ZN(
        vectorData1[52]) );
  AOI22D1BWP U7846 ( .A1(n3576), .A2(\vrf/regTable[5][52] ), .B1(n3567), .B2(
        \vrf/regTable[7][52] ), .ZN(n7314) );
  AOI22D1BWP U7847 ( .A1(n3574), .A2(\vrf/regTable[4][52] ), .B1(n3570), .B2(
        \vrf/regTable[6][52] ), .ZN(n7313) );
  AOI22D1BWP U7848 ( .A1(n3579), .A2(\vrf/regTable[1][52] ), .B1(n3575), .B2(
        \vrf/regTable[3][52] ), .ZN(n7312) );
  AOI22D1BWP U7849 ( .A1(n3581), .A2(\vrf/regTable[0][52] ), .B1(n3572), .B2(
        \vrf/regTable[2][52] ), .ZN(n7311) );
  ND4D1BWP U7850 ( .A1(n7951), .A2(n7952), .A3(n7953), .A4(n7954), .ZN(
        vectorData1[212]) );
  AOI22D1BWP U7851 ( .A1(n3576), .A2(\vrf/regTable[5][212] ), .B1(n3567), .B2(
        \vrf/regTable[7][212] ), .ZN(n7954) );
  AOI22D1BWP U7852 ( .A1(n3574), .A2(\vrf/regTable[4][212] ), .B1(n3570), .B2(
        \vrf/regTable[6][212] ), .ZN(n7953) );
  AOI22D1BWP U7853 ( .A1(n3579), .A2(\vrf/regTable[1][212] ), .B1(n3575), .B2(
        \vrf/regTable[3][212] ), .ZN(n7952) );
  AOI22D1BWP U7854 ( .A1(n3581), .A2(\vrf/regTable[0][212] ), .B1(n3572), .B2(
        \vrf/regTable[2][212] ), .ZN(n7951) );
  ND4D1BWP U7855 ( .A1(n5039), .A2(n5038), .A3(n5037), .A4(n5036), .ZN(n5040)
         );
  AOI22D1BWP U7856 ( .A1(n5185), .A2(vectorData1[84]), .B1(n5230), .B2(
        vectorData1[164]), .ZN(n5036) );
  ND4D1BWP U7857 ( .A1(n7759), .A2(n7760), .A3(n7761), .A4(n7762), .ZN(
        vectorData1[164]) );
  AOI22D1BWP U7858 ( .A1(n3576), .A2(\vrf/regTable[5][164] ), .B1(n3595), .B2(
        \vrf/regTable[7][164] ), .ZN(n7762) );
  AOI22D1BWP U7859 ( .A1(n3574), .A2(\vrf/regTable[4][164] ), .B1(n3596), .B2(
        \vrf/regTable[6][164] ), .ZN(n7761) );
  AOI22D1BWP U7860 ( .A1(n3579), .A2(\vrf/regTable[1][164] ), .B1(n3575), .B2(
        \vrf/regTable[3][164] ), .ZN(n7760) );
  AOI22D1BWP U7861 ( .A1(n3581), .A2(\vrf/regTable[0][164] ), .B1(n3594), .B2(
        \vrf/regTable[2][164] ), .ZN(n7759) );
  ND4D1BWP U7862 ( .A1(n7439), .A2(n7440), .A3(n7441), .A4(n7442), .ZN(
        vectorData1[84]) );
  AOI22D1BWP U7863 ( .A1(n3576), .A2(\vrf/regTable[5][84] ), .B1(n3567), .B2(
        \vrf/regTable[7][84] ), .ZN(n7442) );
  AOI22D1BWP U7864 ( .A1(n3574), .A2(\vrf/regTable[4][84] ), .B1(n3570), .B2(
        \vrf/regTable[6][84] ), .ZN(n7441) );
  AOI22D1BWP U7865 ( .A1(n3579), .A2(\vrf/regTable[1][84] ), .B1(n3575), .B2(
        \vrf/regTable[3][84] ), .ZN(n7440) );
  AOI22D1BWP U7866 ( .A1(n3581), .A2(\vrf/regTable[0][84] ), .B1(n3572), .B2(
        \vrf/regTable[2][84] ), .ZN(n7439) );
  AOI22D1BWP U7867 ( .A1(n5213), .A2(vectorData1[100]), .B1(n5232), .B2(
        vectorData1[148]), .ZN(n5037) );
  ND4D1BWP U7868 ( .A1(n7695), .A2(n7696), .A3(n7697), .A4(n7698), .ZN(
        vectorData1[148]) );
  AOI22D1BWP U7869 ( .A1(n3576), .A2(\vrf/regTable[5][148] ), .B1(n3595), .B2(
        \vrf/regTable[7][148] ), .ZN(n7698) );
  AOI22D1BWP U7870 ( .A1(n3574), .A2(\vrf/regTable[4][148] ), .B1(n3596), .B2(
        \vrf/regTable[6][148] ), .ZN(n7697) );
  AOI22D1BWP U7871 ( .A1(n3579), .A2(\vrf/regTable[1][148] ), .B1(n3599), .B2(
        \vrf/regTable[3][148] ), .ZN(n7696) );
  AOI22D1BWP U7872 ( .A1(n3581), .A2(\vrf/regTable[0][148] ), .B1(n3594), .B2(
        \vrf/regTable[2][148] ), .ZN(n7695) );
  ND4D1BWP U7873 ( .A1(n7503), .A2(n7504), .A3(n7505), .A4(n7506), .ZN(
        vectorData1[100]) );
  AOI22D1BWP U7874 ( .A1(n3576), .A2(\vrf/regTable[5][100] ), .B1(n3595), .B2(
        \vrf/regTable[7][100] ), .ZN(n7506) );
  AOI22D1BWP U7875 ( .A1(n3574), .A2(\vrf/regTable[4][100] ), .B1(n3596), .B2(
        \vrf/regTable[6][100] ), .ZN(n7505) );
  AOI22D1BWP U7876 ( .A1(n3579), .A2(\vrf/regTable[1][100] ), .B1(n3575), .B2(
        \vrf/regTable[3][100] ), .ZN(n7504) );
  AOI22D1BWP U7877 ( .A1(n3581), .A2(\vrf/regTable[0][100] ), .B1(n3594), .B2(
        \vrf/regTable[2][100] ), .ZN(n7503) );
  AOI22D1BWP U7878 ( .A1(n5229), .A2(vectorData1[244]), .B1(n5227), .B2(
        vectorData1[196]), .ZN(n5038) );
  ND4D1BWP U7879 ( .A1(n7887), .A2(n7888), .A3(n7889), .A4(n7890), .ZN(
        vectorData1[196]) );
  AOI22D1BWP U7880 ( .A1(n3576), .A2(\vrf/regTable[5][196] ), .B1(n3595), .B2(
        \vrf/regTable[7][196] ), .ZN(n7890) );
  AOI22D1BWP U7881 ( .A1(n3574), .A2(\vrf/regTable[4][196] ), .B1(n3596), .B2(
        \vrf/regTable[6][196] ), .ZN(n7889) );
  AOI22D1BWP U7882 ( .A1(n3579), .A2(\vrf/regTable[1][196] ), .B1(n3599), .B2(
        \vrf/regTable[3][196] ), .ZN(n7888) );
  AOI22D1BWP U7883 ( .A1(n3581), .A2(\vrf/regTable[0][196] ), .B1(n3594), .B2(
        \vrf/regTable[2][196] ), .ZN(n7887) );
  ND4D1BWP U7884 ( .A1(n8079), .A2(n8080), .A3(n8081), .A4(n8082), .ZN(
        vectorData1[244]) );
  AOI22D1BWP U7885 ( .A1(n3576), .A2(\vrf/regTable[5][244] ), .B1(n3595), .B2(
        \vrf/regTable[7][244] ), .ZN(n8082) );
  AOI22D1BWP U7886 ( .A1(n3574), .A2(\vrf/regTable[4][244] ), .B1(n3596), .B2(
        \vrf/regTable[6][244] ), .ZN(n8081) );
  AOI22D1BWP U7887 ( .A1(n3579), .A2(\vrf/regTable[1][244] ), .B1(n3599), .B2(
        \vrf/regTable[3][244] ), .ZN(n8080) );
  AOI22D1BWP U7888 ( .A1(n3581), .A2(\vrf/regTable[0][244] ), .B1(n3594), .B2(
        \vrf/regTable[2][244] ), .ZN(n8079) );
  AOI22D1BWP U7889 ( .A1(n5226), .A2(vectorData1[132]), .B1(n5233), .B2(
        vectorData1[180]), .ZN(n5039) );
  ND4D1BWP U7890 ( .A1(n7823), .A2(n7824), .A3(n7825), .A4(n7826), .ZN(
        vectorData1[180]) );
  AOI22D1BWP U7891 ( .A1(n3576), .A2(\vrf/regTable[5][180] ), .B1(n3567), .B2(
        \vrf/regTable[7][180] ), .ZN(n7826) );
  AOI22D1BWP U7892 ( .A1(n3574), .A2(\vrf/regTable[4][180] ), .B1(n3570), .B2(
        \vrf/regTable[6][180] ), .ZN(n7825) );
  AOI22D1BWP U7893 ( .A1(n3579), .A2(\vrf/regTable[1][180] ), .B1(n3575), .B2(
        \vrf/regTable[3][180] ), .ZN(n7824) );
  AOI22D1BWP U7894 ( .A1(n3581), .A2(\vrf/regTable[0][180] ), .B1(n3572), .B2(
        \vrf/regTable[2][180] ), .ZN(n7823) );
  ND4D1BWP U7895 ( .A1(n7631), .A2(n7632), .A3(n7633), .A4(n7634), .ZN(
        vectorData1[132]) );
  AOI22D1BWP U7896 ( .A1(n3576), .A2(\vrf/regTable[5][132] ), .B1(n3567), .B2(
        \vrf/regTable[7][132] ), .ZN(n7634) );
  AOI22D1BWP U7897 ( .A1(n3574), .A2(\vrf/regTable[4][132] ), .B1(n3570), .B2(
        \vrf/regTable[6][132] ), .ZN(n7633) );
  AOI22D1BWP U7898 ( .A1(n3579), .A2(\vrf/regTable[1][132] ), .B1(n3599), .B2(
        \vrf/regTable[3][132] ), .ZN(n7632) );
  AOI22D1BWP U7899 ( .A1(n3581), .A2(\vrf/regTable[0][132] ), .B1(n3572), .B2(
        \vrf/regTable[2][132] ), .ZN(n7631) );
  ND4D1BWP U7900 ( .A1(n7247), .A2(n7248), .A3(n7249), .A4(n7250), .ZN(
        vectorData1[36]) );
  AOI22D1BWP U7901 ( .A1(n3576), .A2(\vrf/regTable[5][36] ), .B1(n3567), .B2(
        \vrf/regTable[7][36] ), .ZN(n7250) );
  AOI22D1BWP U7902 ( .A1(n3574), .A2(\vrf/regTable[4][36] ), .B1(n3570), .B2(
        \vrf/regTable[6][36] ), .ZN(n7249) );
  AOI22D1BWP U7903 ( .A1(n3579), .A2(\vrf/regTable[1][36] ), .B1(n3575), .B2(
        \vrf/regTable[3][36] ), .ZN(n7248) );
  AOI22D1BWP U7904 ( .A1(n3581), .A2(\vrf/regTable[0][36] ), .B1(n3572), .B2(
        \vrf/regTable[2][36] ), .ZN(n7247) );
  AOI22D1BWP U7905 ( .A1(n5231), .A2(vectorData1[116]), .B1(n5184), .B2(
        vectorData1[20]), .ZN(n5041) );
  ND4D1BWP U7906 ( .A1(n7183), .A2(n7184), .A3(n7185), .A4(n7186), .ZN(
        vectorData1[20]) );
  AOI22D1BWP U7907 ( .A1(n3576), .A2(\vrf/regTable[5][20] ), .B1(n3567), .B2(
        \vrf/regTable[7][20] ), .ZN(n7186) );
  AOI22D1BWP U7908 ( .A1(n3574), .A2(\vrf/regTable[4][20] ), .B1(n3570), .B2(
        \vrf/regTable[6][20] ), .ZN(n7185) );
  AOI22D1BWP U7909 ( .A1(n3579), .A2(\vrf/regTable[1][20] ), .B1(n3575), .B2(
        \vrf/regTable[3][20] ), .ZN(n7184) );
  AOI22D1BWP U7910 ( .A1(n3581), .A2(\vrf/regTable[0][20] ), .B1(n3572), .B2(
        \vrf/regTable[2][20] ), .ZN(n7183) );
  ND4D1BWP U7911 ( .A1(n7567), .A2(n7568), .A3(n7569), .A4(n7570), .ZN(
        vectorData1[116]) );
  AOI22D1BWP U7912 ( .A1(n3576), .A2(\vrf/regTable[5][116] ), .B1(n3595), .B2(
        \vrf/regTable[7][116] ), .ZN(n7570) );
  AOI22D1BWP U7913 ( .A1(n3574), .A2(\vrf/regTable[4][116] ), .B1(n3596), .B2(
        \vrf/regTable[6][116] ), .ZN(n7569) );
  AOI22D1BWP U7914 ( .A1(n3579), .A2(\vrf/regTable[1][116] ), .B1(n3599), .B2(
        \vrf/regTable[3][116] ), .ZN(n7568) );
  AOI22D1BWP U7915 ( .A1(n3581), .A2(\vrf/regTable[0][116] ), .B1(n3594), .B2(
        \vrf/regTable[2][116] ), .ZN(n7567) );
  ND4D1BWP U7916 ( .A1(n8015), .A2(n8016), .A3(n8017), .A4(n8018), .ZN(
        vectorData1[228]) );
  AOI22D1BWP U7917 ( .A1(n3576), .A2(\vrf/regTable[5][228] ), .B1(n3595), .B2(
        \vrf/regTable[7][228] ), .ZN(n8018) );
  AOI22D1BWP U7918 ( .A1(n3574), .A2(\vrf/regTable[4][228] ), .B1(n3596), .B2(
        \vrf/regTable[6][228] ), .ZN(n8017) );
  AOI22D1BWP U7919 ( .A1(n3579), .A2(\vrf/regTable[1][228] ), .B1(n3599), .B2(
        \vrf/regTable[3][228] ), .ZN(n8016) );
  AOI22D1BWP U7920 ( .A1(n3581), .A2(\vrf/regTable[0][228] ), .B1(n3594), .B2(
        \vrf/regTable[2][228] ), .ZN(n8015) );
  AO222D1BWP U7921 ( .A1(n3641), .A2(n4548), .B1(n5527), .B2(n4628), .C1(n3669), .C2(vectorToLoad[103]), .Z(N4320) );
  NR2XD0BWP U7922 ( .A1(n4655), .A2(n5282), .ZN(n5527) );
  OAI211D1BWP U7923 ( .A1(n5350), .A2(n5509), .B(n5351), .C(n4406), .ZN(N4370)
         );
  AOI22D1BWP U7924 ( .A1(n3669), .A2(vectorToLoad[152]), .B1(n4626), .B2(n5400), .ZN(n5351) );
  NR2XD0BWP U7925 ( .A1(n5275), .A2(cycles[0]), .ZN(n5400) );
  AO211D1BWP U7926 ( .A1(n4073), .A2(scalarData1[3]), .B(n3825), .C(n3824), 
        .Z(N4179) );
  MOAI22D0BWP U7927 ( .A1(n3830), .A2(n3823), .B1(n4072), .B2(vectorData1[3]), 
        .ZN(n3824) );
  ND4D1BWP U7928 ( .A1(n7131), .A2(n7132), .A3(n7133), .A4(n7134), .ZN(
        vectorData1[3]) );
  AOI22D1BWP U7929 ( .A1(n3576), .A2(\vrf/regTable[5][3] ), .B1(n3595), .B2(
        \vrf/regTable[7][3] ), .ZN(n7134) );
  AOI22D1BWP U7930 ( .A1(n3574), .A2(\vrf/regTable[4][3] ), .B1(n3596), .B2(
        \vrf/regTable[6][3] ), .ZN(n7133) );
  AOI22D1BWP U7931 ( .A1(n3579), .A2(\vrf/regTable[1][3] ), .B1(n3599), .B2(
        \vrf/regTable[3][3] ), .ZN(n7132) );
  AOI22D1BWP U7932 ( .A1(n3581), .A2(\vrf/regTable[0][3] ), .B1(n3594), .B2(
        \vrf/regTable[2][3] ), .ZN(n7131) );
  AOI31D1BWP U7933 ( .A1(n5034), .A2(n5033), .A3(n5035), .B(n4070), .ZN(n3825)
         );
  AOI22D1BWP U7934 ( .A1(n5230), .A2(vectorData1[163]), .B1(n5186), .B2(
        vectorData1[67]), .ZN(n5035) );
  ND4D1BWP U7935 ( .A1(n7371), .A2(n7372), .A3(n7373), .A4(n7374), .ZN(
        vectorData1[67]) );
  AOI22D1BWP U7936 ( .A1(n3576), .A2(\vrf/regTable[5][67] ), .B1(n3595), .B2(
        \vrf/regTable[7][67] ), .ZN(n7374) );
  AOI22D1BWP U7937 ( .A1(n3574), .A2(\vrf/regTable[4][67] ), .B1(n3596), .B2(
        \vrf/regTable[6][67] ), .ZN(n7373) );
  AOI22D1BWP U7938 ( .A1(n3579), .A2(\vrf/regTable[1][67] ), .B1(n3599), .B2(
        \vrf/regTable[3][67] ), .ZN(n7372) );
  AOI22D1BWP U7939 ( .A1(n3581), .A2(\vrf/regTable[0][67] ), .B1(n3594), .B2(
        \vrf/regTable[2][67] ), .ZN(n7371) );
  ND4D1BWP U7940 ( .A1(n7755), .A2(n7756), .A3(n7757), .A4(n7758), .ZN(
        vectorData1[163]) );
  AOI22D1BWP U7941 ( .A1(n3576), .A2(\vrf/regTable[5][163] ), .B1(n3595), .B2(
        \vrf/regTable[7][163] ), .ZN(n7758) );
  AOI22D1BWP U7942 ( .A1(n3574), .A2(\vrf/regTable[4][163] ), .B1(n3596), .B2(
        \vrf/regTable[6][163] ), .ZN(n7757) );
  AOI22D1BWP U7943 ( .A1(n3579), .A2(\vrf/regTable[1][163] ), .B1(n3575), .B2(
        \vrf/regTable[3][163] ), .ZN(n7756) );
  AOI22D1BWP U7944 ( .A1(n3581), .A2(\vrf/regTable[0][163] ), .B1(n3594), .B2(
        \vrf/regTable[2][163] ), .ZN(n7755) );
  AOI211XD0BWP U7945 ( .A1(n5213), .A2(vectorData1[99]), .B(n5032), .C(n5031), 
        .ZN(n5033) );
  ND4D1BWP U7946 ( .A1(n5030), .A2(n5029), .A3(n5028), .A4(n5027), .ZN(n5031)
         );
  AOI22D1BWP U7947 ( .A1(n5226), .A2(vectorData1[131]), .B1(n5185), .B2(
        vectorData1[83]), .ZN(n5027) );
  ND4D1BWP U7948 ( .A1(n7435), .A2(n7436), .A3(n7437), .A4(n7438), .ZN(
        vectorData1[83]) );
  AOI22D1BWP U7949 ( .A1(n3576), .A2(\vrf/regTable[5][83] ), .B1(n3595), .B2(
        \vrf/regTable[7][83] ), .ZN(n7438) );
  AOI22D1BWP U7950 ( .A1(n3574), .A2(\vrf/regTable[4][83] ), .B1(n3596), .B2(
        \vrf/regTable[6][83] ), .ZN(n7437) );
  AOI22D1BWP U7951 ( .A1(n3579), .A2(\vrf/regTable[1][83] ), .B1(n3599), .B2(
        \vrf/regTable[3][83] ), .ZN(n7436) );
  AOI22D1BWP U7952 ( .A1(n3581), .A2(\vrf/regTable[0][83] ), .B1(n3594), .B2(
        \vrf/regTable[2][83] ), .ZN(n7435) );
  ND4D1BWP U7953 ( .A1(n7627), .A2(n7628), .A3(n7629), .A4(n7630), .ZN(
        vectorData1[131]) );
  AOI22D1BWP U7954 ( .A1(n3576), .A2(\vrf/regTable[5][131] ), .B1(n3567), .B2(
        \vrf/regTable[7][131] ), .ZN(n7630) );
  AOI22D1BWP U7955 ( .A1(n3574), .A2(\vrf/regTable[4][131] ), .B1(n3570), .B2(
        \vrf/regTable[6][131] ), .ZN(n7629) );
  AOI22D1BWP U7956 ( .A1(n3579), .A2(\vrf/regTable[1][131] ), .B1(n3575), .B2(
        \vrf/regTable[3][131] ), .ZN(n7628) );
  AOI22D1BWP U7957 ( .A1(n3581), .A2(\vrf/regTable[0][131] ), .B1(n3572), .B2(
        \vrf/regTable[2][131] ), .ZN(n7627) );
  AOI22D1BWP U7958 ( .A1(n5188), .A2(vectorData1[51]), .B1(n5227), .B2(
        vectorData1[195]), .ZN(n5028) );
  ND4D1BWP U7959 ( .A1(n7883), .A2(n7884), .A3(n7885), .A4(n7886), .ZN(
        vectorData1[195]) );
  AOI22D1BWP U7960 ( .A1(n3576), .A2(\vrf/regTable[5][195] ), .B1(n3595), .B2(
        \vrf/regTable[7][195] ), .ZN(n7886) );
  AOI22D1BWP U7961 ( .A1(n3574), .A2(\vrf/regTable[4][195] ), .B1(n3596), .B2(
        \vrf/regTable[6][195] ), .ZN(n7885) );
  AOI22D1BWP U7962 ( .A1(n3579), .A2(\vrf/regTable[1][195] ), .B1(n3599), .B2(
        \vrf/regTable[3][195] ), .ZN(n7884) );
  AOI22D1BWP U7963 ( .A1(n3581), .A2(\vrf/regTable[0][195] ), .B1(n3594), .B2(
        \vrf/regTable[2][195] ), .ZN(n7883) );
  ND4D1BWP U7964 ( .A1(n7307), .A2(n7308), .A3(n7309), .A4(n7310), .ZN(
        vectorData1[51]) );
  AOI22D1BWP U7965 ( .A1(n3576), .A2(\vrf/regTable[5][51] ), .B1(n3595), .B2(
        \vrf/regTable[7][51] ), .ZN(n7310) );
  AOI22D1BWP U7966 ( .A1(n3574), .A2(\vrf/regTable[4][51] ), .B1(n3596), .B2(
        \vrf/regTable[6][51] ), .ZN(n7309) );
  AOI22D1BWP U7967 ( .A1(n3579), .A2(\vrf/regTable[1][51] ), .B1(n3599), .B2(
        \vrf/regTable[3][51] ), .ZN(n7308) );
  AOI22D1BWP U7968 ( .A1(n3581), .A2(\vrf/regTable[0][51] ), .B1(n3594), .B2(
        \vrf/regTable[2][51] ), .ZN(n7307) );
  AOI22D1BWP U7969 ( .A1(n5228), .A2(vectorData1[211]), .B1(n3601), .B2(
        vectorData1[35]), .ZN(n5029) );
  ND4D1BWP U7970 ( .A1(n7243), .A2(n7244), .A3(n7245), .A4(n7246), .ZN(
        vectorData1[35]) );
  AOI22D1BWP U7971 ( .A1(n3576), .A2(\vrf/regTable[5][35] ), .B1(n3567), .B2(
        \vrf/regTable[7][35] ), .ZN(n7246) );
  AOI22D1BWP U7972 ( .A1(n3574), .A2(\vrf/regTable[4][35] ), .B1(n3570), .B2(
        \vrf/regTable[6][35] ), .ZN(n7245) );
  AOI22D1BWP U7973 ( .A1(n3579), .A2(\vrf/regTable[1][35] ), .B1(n3575), .B2(
        \vrf/regTable[3][35] ), .ZN(n7244) );
  AOI22D1BWP U7974 ( .A1(n3581), .A2(\vrf/regTable[0][35] ), .B1(n3572), .B2(
        \vrf/regTable[2][35] ), .ZN(n7243) );
  ND4D1BWP U7975 ( .A1(n7947), .A2(n7948), .A3(n7949), .A4(n7950), .ZN(
        vectorData1[211]) );
  AOI22D1BWP U7976 ( .A1(n3576), .A2(\vrf/regTable[5][211] ), .B1(n7118), .B2(
        \vrf/regTable[7][211] ), .ZN(n7950) );
  AOI22D1BWP U7977 ( .A1(n3574), .A2(\vrf/regTable[4][211] ), .B1(n7116), .B2(
        \vrf/regTable[6][211] ), .ZN(n7949) );
  AOI22D1BWP U7978 ( .A1(n3579), .A2(\vrf/regTable[1][211] ), .B1(n7114), .B2(
        \vrf/regTable[3][211] ), .ZN(n7948) );
  AOI22D1BWP U7979 ( .A1(n3581), .A2(\vrf/regTable[0][211] ), .B1(n7110), .B2(
        \vrf/regTable[2][211] ), .ZN(n7947) );
  AOI22D1BWP U7980 ( .A1(n5231), .A2(vectorData1[115]), .B1(n5233), .B2(
        vectorData1[179]), .ZN(n5030) );
  ND4D1BWP U7981 ( .A1(n7819), .A2(n7820), .A3(n7821), .A4(n7822), .ZN(
        vectorData1[179]) );
  AOI22D1BWP U7982 ( .A1(n3576), .A2(\vrf/regTable[5][179] ), .B1(n3595), .B2(
        \vrf/regTable[7][179] ), .ZN(n7822) );
  AOI22D1BWP U7983 ( .A1(n3574), .A2(\vrf/regTable[4][179] ), .B1(n3596), .B2(
        \vrf/regTable[6][179] ), .ZN(n7821) );
  AOI22D1BWP U7984 ( .A1(n3579), .A2(\vrf/regTable[1][179] ), .B1(n3599), .B2(
        \vrf/regTable[3][179] ), .ZN(n7820) );
  AOI22D1BWP U7985 ( .A1(n3581), .A2(\vrf/regTable[0][179] ), .B1(n3594), .B2(
        \vrf/regTable[2][179] ), .ZN(n7819) );
  ND4D1BWP U7986 ( .A1(n7563), .A2(n7564), .A3(n7565), .A4(n7566), .ZN(
        vectorData1[115]) );
  AOI22D1BWP U7987 ( .A1(n3576), .A2(\vrf/regTable[5][115] ), .B1(n3567), .B2(
        \vrf/regTable[7][115] ), .ZN(n7566) );
  AOI22D1BWP U7988 ( .A1(n3574), .A2(\vrf/regTable[4][115] ), .B1(n3570), .B2(
        \vrf/regTable[6][115] ), .ZN(n7565) );
  AOI22D1BWP U7989 ( .A1(n3579), .A2(\vrf/regTable[1][115] ), .B1(n3599), .B2(
        \vrf/regTable[3][115] ), .ZN(n7564) );
  AOI22D1BWP U7990 ( .A1(n3581), .A2(\vrf/regTable[0][115] ), .B1(n3572), .B2(
        \vrf/regTable[2][115] ), .ZN(n7563) );
  AO22D1BWP U7991 ( .A1(n5184), .A2(vectorData1[19]), .B1(n5232), .B2(
        vectorData1[147]), .Z(n5032) );
  ND4D1BWP U7992 ( .A1(n7691), .A2(n7692), .A3(n7693), .A4(n7694), .ZN(
        vectorData1[147]) );
  AOI22D1BWP U7993 ( .A1(n3576), .A2(\vrf/regTable[5][147] ), .B1(n3595), .B2(
        \vrf/regTable[7][147] ), .ZN(n7694) );
  AOI22D1BWP U7994 ( .A1(n3574), .A2(\vrf/regTable[4][147] ), .B1(n3596), .B2(
        \vrf/regTable[6][147] ), .ZN(n7693) );
  AOI22D1BWP U7995 ( .A1(n3579), .A2(\vrf/regTable[1][147] ), .B1(n3599), .B2(
        \vrf/regTable[3][147] ), .ZN(n7692) );
  AOI22D1BWP U7996 ( .A1(n3581), .A2(\vrf/regTable[0][147] ), .B1(n3594), .B2(
        \vrf/regTable[2][147] ), .ZN(n7691) );
  ND4D1BWP U7997 ( .A1(n7179), .A2(n7180), .A3(n7181), .A4(n7182), .ZN(
        vectorData1[19]) );
  AOI22D1BWP U7998 ( .A1(n7117), .A2(\vrf/regTable[5][19] ), .B1(n3595), .B2(
        \vrf/regTable[7][19] ), .ZN(n7182) );
  AOI22D1BWP U7999 ( .A1(n3574), .A2(\vrf/regTable[4][19] ), .B1(n3596), .B2(
        \vrf/regTable[6][19] ), .ZN(n7181) );
  AOI22D1BWP U8000 ( .A1(n7112), .A2(\vrf/regTable[1][19] ), .B1(n3599), .B2(
        \vrf/regTable[3][19] ), .ZN(n7180) );
  AOI22D1BWP U8001 ( .A1(n3581), .A2(\vrf/regTable[0][19] ), .B1(n3594), .B2(
        \vrf/regTable[2][19] ), .ZN(n7179) );
  ND4D1BWP U8002 ( .A1(n7499), .A2(n7500), .A3(n7501), .A4(n7502), .ZN(
        vectorData1[99]) );
  AOI22D1BWP U8003 ( .A1(n3576), .A2(\vrf/regTable[5][99] ), .B1(n3567), .B2(
        \vrf/regTable[7][99] ), .ZN(n7502) );
  AOI22D1BWP U8004 ( .A1(n3574), .A2(\vrf/regTable[4][99] ), .B1(n3570), .B2(
        \vrf/regTable[6][99] ), .ZN(n7501) );
  AOI22D1BWP U8005 ( .A1(n3579), .A2(\vrf/regTable[1][99] ), .B1(n3575), .B2(
        \vrf/regTable[3][99] ), .ZN(n7500) );
  AOI22D1BWP U8006 ( .A1(n3581), .A2(\vrf/regTable[0][99] ), .B1(n3572), .B2(
        \vrf/regTable[2][99] ), .ZN(n7499) );
  AOI22D1BWP U8007 ( .A1(n5229), .A2(vectorData1[243]), .B1(n5187), .B2(
        vectorData1[227]), .ZN(n5034) );
  ND4D1BWP U8008 ( .A1(n8011), .A2(n8012), .A3(n8013), .A4(n8014), .ZN(
        vectorData1[227]) );
  AOI22D1BWP U8009 ( .A1(n3576), .A2(\vrf/regTable[5][227] ), .B1(n3567), .B2(
        \vrf/regTable[7][227] ), .ZN(n8014) );
  AOI22D1BWP U8010 ( .A1(n3574), .A2(\vrf/regTable[4][227] ), .B1(n3570), .B2(
        \vrf/regTable[6][227] ), .ZN(n8013) );
  AOI22D1BWP U8011 ( .A1(n3579), .A2(\vrf/regTable[1][227] ), .B1(n3575), .B2(
        \vrf/regTable[3][227] ), .ZN(n8012) );
  AOI22D1BWP U8012 ( .A1(n3581), .A2(\vrf/regTable[0][227] ), .B1(n3572), .B2(
        \vrf/regTable[2][227] ), .ZN(n8011) );
  ND4D1BWP U8013 ( .A1(n8075), .A2(n8076), .A3(n8077), .A4(n8078), .ZN(
        vectorData1[243]) );
  AOI22D1BWP U8014 ( .A1(n3576), .A2(\vrf/regTable[5][243] ), .B1(n3567), .B2(
        \vrf/regTable[7][243] ), .ZN(n8078) );
  AOI22D1BWP U8015 ( .A1(n3574), .A2(\vrf/regTable[4][243] ), .B1(n3570), .B2(
        \vrf/regTable[6][243] ), .ZN(n8077) );
  AOI22D1BWP U8016 ( .A1(n3579), .A2(\vrf/regTable[1][243] ), .B1(n3575), .B2(
        \vrf/regTable[3][243] ), .ZN(n8076) );
  AOI22D1BWP U8017 ( .A1(n3581), .A2(\vrf/regTable[0][243] ), .B1(n3572), .B2(
        \vrf/regTable[2][243] ), .ZN(n8075) );
  ND4D1BWP U8018 ( .A1(n8301), .A2(n8302), .A3(n8303), .A4(n8304), .ZN(
        scalarData1[3]) );
  AOI22D1BWP U8019 ( .A1(n8287), .A2(\srf/regTable[5][3] ), .B1(n8288), .B2(
        \srf/regTable[7][3] ), .ZN(n8304) );
  AOI22D1BWP U8020 ( .A1(n8285), .A2(\srf/regTable[4][3] ), .B1(n8286), .B2(
        \srf/regTable[6][3] ), .ZN(n8303) );
  AOI22D1BWP U8021 ( .A1(n8282), .A2(\srf/regTable[1][3] ), .B1(n8284), .B2(
        \srf/regTable[3][3] ), .ZN(n8302) );
  AOI22D1BWP U8022 ( .A1(n8278), .A2(\srf/regTable[0][3] ), .B1(n8280), .B2(
        \srf/regTable[2][3] ), .ZN(n8301) );
  OAI211D1BWP U8023 ( .A1(n5491), .A2(n4405), .B(n5354), .C(n4535), .ZN(N4371)
         );
  AOI22D1BWP U8024 ( .A1(n3669), .A2(vectorToLoad[153]), .B1(n4627), .B2(n5353), .ZN(n5354) );
  NR2XD0BWP U8025 ( .A1(n5334), .A2(n4651), .ZN(n5353) );
  NR2XD0BWP U8026 ( .A1(n5276), .A2(cycles[0]), .ZN(n5352) );
  AO222D1BWP U8027 ( .A1(n3669), .A2(vectorToLoad[48]), .B1(n5289), .B2(n3649), 
        .C1(n4549), .C2(n5536), .Z(N4265) );
  AOI21D1BWP U8028 ( .A1(cycles[1]), .A2(n5284), .B(n136), .ZN(n5536) );
  AOI21D1BWP U8029 ( .A1(n4642), .A2(n137), .B(n5253), .ZN(n5284) );
  NR2XD0BWP U8030 ( .A1(n6004), .A2(n3679), .ZN(n5253) );
  OAI211D1BWP U8031 ( .A1(n5355), .A2(n5509), .B(n5356), .C(n4406), .ZN(N4372)
         );
  AOI22D1BWP U8032 ( .A1(n3668), .A2(vectorToLoad[154]), .B1(n4626), .B2(n5403), .ZN(n5356) );
  NR2XD0BWP U8033 ( .A1(n5277), .A2(cycles[0]), .ZN(n5403) );
  AO211D1BWP U8034 ( .A1(n4073), .A2(scalarData1[2]), .B(n3810), .C(n3809), 
        .Z(N4178) );
  MOAI22D0BWP U8035 ( .A1(n3830), .A2(n3808), .B1(n4072), .B2(vectorData1[2]), 
        .ZN(n3809) );
  ND4D1BWP U8036 ( .A1(n7127), .A2(n7128), .A3(n7129), .A4(n7130), .ZN(
        vectorData1[2]) );
  AOI22D1BWP U8037 ( .A1(n3576), .A2(\vrf/regTable[5][2] ), .B1(n3595), .B2(
        \vrf/regTable[7][2] ), .ZN(n7130) );
  AOI22D1BWP U8038 ( .A1(n3574), .A2(\vrf/regTable[4][2] ), .B1(n3596), .B2(
        \vrf/regTable[6][2] ), .ZN(n7129) );
  AOI22D1BWP U8039 ( .A1(n3579), .A2(\vrf/regTable[1][2] ), .B1(n3599), .B2(
        \vrf/regTable[3][2] ), .ZN(n7128) );
  AOI22D1BWP U8040 ( .A1(n3581), .A2(\vrf/regTable[0][2] ), .B1(n3594), .B2(
        \vrf/regTable[2][2] ), .ZN(n7127) );
  AOI31D1BWP U8041 ( .A1(n5025), .A2(n5024), .A3(n5026), .B(n4070), .ZN(n3810)
         );
  AOI22D1BWP U8042 ( .A1(n5213), .A2(vectorData1[98]), .B1(n5232), .B2(
        vectorData1[146]), .ZN(n5026) );
  ND4D1BWP U8043 ( .A1(n7687), .A2(n7688), .A3(n7689), .A4(n7690), .ZN(
        vectorData1[146]) );
  AOI22D1BWP U8044 ( .A1(n3576), .A2(\vrf/regTable[5][146] ), .B1(n3595), .B2(
        \vrf/regTable[7][146] ), .ZN(n7690) );
  AOI22D1BWP U8045 ( .A1(n3574), .A2(\vrf/regTable[4][146] ), .B1(n3596), .B2(
        \vrf/regTable[6][146] ), .ZN(n7689) );
  AOI22D1BWP U8046 ( .A1(n3579), .A2(\vrf/regTable[1][146] ), .B1(n3599), .B2(
        \vrf/regTable[3][146] ), .ZN(n7688) );
  AOI22D1BWP U8047 ( .A1(n3581), .A2(\vrf/regTable[0][146] ), .B1(n3594), .B2(
        \vrf/regTable[2][146] ), .ZN(n7687) );
  ND4D1BWP U8048 ( .A1(n7495), .A2(n7496), .A3(n7497), .A4(n7498), .ZN(
        vectorData1[98]) );
  AOI22D1BWP U8049 ( .A1(n3576), .A2(\vrf/regTable[5][98] ), .B1(n3567), .B2(
        \vrf/regTable[7][98] ), .ZN(n7498) );
  AOI22D1BWP U8050 ( .A1(n3574), .A2(\vrf/regTable[4][98] ), .B1(n3570), .B2(
        \vrf/regTable[6][98] ), .ZN(n7497) );
  AOI22D1BWP U8051 ( .A1(n3579), .A2(\vrf/regTable[1][98] ), .B1(n3575), .B2(
        \vrf/regTable[3][98] ), .ZN(n7496) );
  AOI22D1BWP U8052 ( .A1(n3581), .A2(\vrf/regTable[0][98] ), .B1(n3572), .B2(
        \vrf/regTable[2][98] ), .ZN(n7495) );
  AOI211XD0BWP U8053 ( .A1(n5229), .A2(vectorData1[242]), .B(n5023), .C(n5022), 
        .ZN(n5024) );
  ND4D1BWP U8054 ( .A1(n5021), .A2(n5020), .A3(n5019), .A4(n5018), .ZN(n5022)
         );
  AOI22D1BWP U8055 ( .A1(n5228), .A2(vectorData1[210]), .B1(n5230), .B2(
        vectorData1[162]), .ZN(n5018) );
  ND4D1BWP U8056 ( .A1(n7751), .A2(n7752), .A3(n7753), .A4(n7754), .ZN(
        vectorData1[162]) );
  AOI22D1BWP U8057 ( .A1(n3576), .A2(\vrf/regTable[5][162] ), .B1(n3567), .B2(
        \vrf/regTable[7][162] ), .ZN(n7754) );
  AOI22D1BWP U8058 ( .A1(n3574), .A2(\vrf/regTable[4][162] ), .B1(n3570), .B2(
        \vrf/regTable[6][162] ), .ZN(n7753) );
  AOI22D1BWP U8059 ( .A1(n3579), .A2(\vrf/regTable[1][162] ), .B1(n3575), .B2(
        \vrf/regTable[3][162] ), .ZN(n7752) );
  AOI22D1BWP U8060 ( .A1(n3581), .A2(\vrf/regTable[0][162] ), .B1(n3572), .B2(
        \vrf/regTable[2][162] ), .ZN(n7751) );
  ND4D1BWP U8061 ( .A1(n7943), .A2(n7944), .A3(n7945), .A4(n7946), .ZN(
        vectorData1[210]) );
  AOI22D1BWP U8062 ( .A1(n3576), .A2(\vrf/regTable[5][210] ), .B1(n7118), .B2(
        \vrf/regTable[7][210] ), .ZN(n7946) );
  AOI22D1BWP U8063 ( .A1(n3574), .A2(\vrf/regTable[4][210] ), .B1(n7116), .B2(
        \vrf/regTable[6][210] ), .ZN(n7945) );
  AOI22D1BWP U8064 ( .A1(n3579), .A2(\vrf/regTable[1][210] ), .B1(n7114), .B2(
        \vrf/regTable[3][210] ), .ZN(n7944) );
  AOI22D1BWP U8065 ( .A1(n3581), .A2(\vrf/regTable[0][210] ), .B1(n7110), .B2(
        \vrf/regTable[2][210] ), .ZN(n7943) );
  AOI22D1BWP U8066 ( .A1(n5226), .A2(vectorData1[130]), .B1(n3601), .B2(
        vectorData1[34]), .ZN(n5019) );
  ND4D1BWP U8067 ( .A1(n7239), .A2(n7240), .A3(n7241), .A4(n7242), .ZN(
        vectorData1[34]) );
  AOI22D1BWP U8068 ( .A1(n3576), .A2(\vrf/regTable[5][34] ), .B1(n3595), .B2(
        \vrf/regTable[7][34] ), .ZN(n7242) );
  AOI22D1BWP U8069 ( .A1(n3574), .A2(\vrf/regTable[4][34] ), .B1(n3596), .B2(
        \vrf/regTable[6][34] ), .ZN(n7241) );
  AOI22D1BWP U8070 ( .A1(n3579), .A2(\vrf/regTable[1][34] ), .B1(n3599), .B2(
        \vrf/regTable[3][34] ), .ZN(n7240) );
  AOI22D1BWP U8071 ( .A1(n3581), .A2(\vrf/regTable[0][34] ), .B1(n3594), .B2(
        \vrf/regTable[2][34] ), .ZN(n7239) );
  ND4D1BWP U8072 ( .A1(n7623), .A2(n7624), .A3(n7625), .A4(n7626), .ZN(
        vectorData1[130]) );
  AOI22D1BWP U8073 ( .A1(n3576), .A2(\vrf/regTable[5][130] ), .B1(n3567), .B2(
        \vrf/regTable[7][130] ), .ZN(n7626) );
  AOI22D1BWP U8074 ( .A1(n3574), .A2(\vrf/regTable[4][130] ), .B1(n3570), .B2(
        \vrf/regTable[6][130] ), .ZN(n7625) );
  AOI22D1BWP U8075 ( .A1(n3579), .A2(\vrf/regTable[1][130] ), .B1(n3575), .B2(
        \vrf/regTable[3][130] ), .ZN(n7624) );
  AOI22D1BWP U8076 ( .A1(n3581), .A2(\vrf/regTable[0][130] ), .B1(n3572), .B2(
        \vrf/regTable[2][130] ), .ZN(n7623) );
  AOI22D1BWP U8077 ( .A1(n5185), .A2(vectorData1[82]), .B1(n5233), .B2(
        vectorData1[178]), .ZN(n5020) );
  ND4D1BWP U8078 ( .A1(n7815), .A2(n7816), .A3(n7817), .A4(n7818), .ZN(
        vectorData1[178]) );
  AOI22D1BWP U8079 ( .A1(n3576), .A2(\vrf/regTable[5][178] ), .B1(n3595), .B2(
        \vrf/regTable[7][178] ), .ZN(n7818) );
  AOI22D1BWP U8080 ( .A1(n3574), .A2(\vrf/regTable[4][178] ), .B1(n3596), .B2(
        \vrf/regTable[6][178] ), .ZN(n7817) );
  AOI22D1BWP U8081 ( .A1(n3579), .A2(\vrf/regTable[1][178] ), .B1(n3599), .B2(
        \vrf/regTable[3][178] ), .ZN(n7816) );
  AOI22D1BWP U8082 ( .A1(n3581), .A2(\vrf/regTable[0][178] ), .B1(n3594), .B2(
        \vrf/regTable[2][178] ), .ZN(n7815) );
  ND4D1BWP U8083 ( .A1(n7431), .A2(n7432), .A3(n7433), .A4(n7434), .ZN(
        vectorData1[82]) );
  AOI22D1BWP U8084 ( .A1(n7117), .A2(\vrf/regTable[5][82] ), .B1(n3567), .B2(
        \vrf/regTable[7][82] ), .ZN(n7434) );
  AOI22D1BWP U8085 ( .A1(n7115), .A2(\vrf/regTable[4][82] ), .B1(n3570), .B2(
        \vrf/regTable[6][82] ), .ZN(n7433) );
  AOI22D1BWP U8086 ( .A1(n7112), .A2(\vrf/regTable[1][82] ), .B1(n3575), .B2(
        \vrf/regTable[3][82] ), .ZN(n7432) );
  AOI22D1BWP U8087 ( .A1(n7108), .A2(\vrf/regTable[0][82] ), .B1(n3572), .B2(
        \vrf/regTable[2][82] ), .ZN(n7431) );
  AOI22D1BWP U8088 ( .A1(n5187), .A2(vectorData1[226]), .B1(n5186), .B2(
        vectorData1[66]), .ZN(n5021) );
  ND4D1BWP U8089 ( .A1(n7367), .A2(n7368), .A3(n7369), .A4(n7370), .ZN(
        vectorData1[66]) );
  AOI22D1BWP U8090 ( .A1(n7117), .A2(\vrf/regTable[5][66] ), .B1(n3567), .B2(
        \vrf/regTable[7][66] ), .ZN(n7370) );
  AOI22D1BWP U8091 ( .A1(n7115), .A2(\vrf/regTable[4][66] ), .B1(n3570), .B2(
        \vrf/regTable[6][66] ), .ZN(n7369) );
  AOI22D1BWP U8092 ( .A1(n7112), .A2(\vrf/regTable[1][66] ), .B1(n3575), .B2(
        \vrf/regTable[3][66] ), .ZN(n7368) );
  AOI22D1BWP U8093 ( .A1(n7108), .A2(\vrf/regTable[0][66] ), .B1(n3572), .B2(
        \vrf/regTable[2][66] ), .ZN(n7367) );
  ND4D1BWP U8094 ( .A1(n8007), .A2(n8008), .A3(n8009), .A4(n8010), .ZN(
        vectorData1[226]) );
  AOI22D1BWP U8095 ( .A1(n3576), .A2(\vrf/regTable[5][226] ), .B1(n3567), .B2(
        \vrf/regTable[7][226] ), .ZN(n8010) );
  AOI22D1BWP U8096 ( .A1(n3574), .A2(\vrf/regTable[4][226] ), .B1(n3570), .B2(
        \vrf/regTable[6][226] ), .ZN(n8009) );
  AOI22D1BWP U8097 ( .A1(n3579), .A2(\vrf/regTable[1][226] ), .B1(n3575), .B2(
        \vrf/regTable[3][226] ), .ZN(n8008) );
  AOI22D1BWP U8098 ( .A1(n3581), .A2(\vrf/regTable[0][226] ), .B1(n3572), .B2(
        \vrf/regTable[2][226] ), .ZN(n8007) );
  AO22D1BWP U8099 ( .A1(n5188), .A2(vectorData1[50]), .B1(n5227), .B2(
        vectorData1[194]), .Z(n5023) );
  ND4D1BWP U8100 ( .A1(n7879), .A2(n7880), .A3(n7881), .A4(n7882), .ZN(
        vectorData1[194]) );
  AOI22D1BWP U8101 ( .A1(n3576), .A2(\vrf/regTable[5][194] ), .B1(n3567), .B2(
        \vrf/regTable[7][194] ), .ZN(n7882) );
  AOI22D1BWP U8102 ( .A1(n3574), .A2(\vrf/regTable[4][194] ), .B1(n3570), .B2(
        \vrf/regTable[6][194] ), .ZN(n7881) );
  AOI22D1BWP U8103 ( .A1(n3579), .A2(\vrf/regTable[1][194] ), .B1(n3575), .B2(
        \vrf/regTable[3][194] ), .ZN(n7880) );
  AOI22D1BWP U8104 ( .A1(n3581), .A2(\vrf/regTable[0][194] ), .B1(n3572), .B2(
        \vrf/regTable[2][194] ), .ZN(n7879) );
  ND4D1BWP U8105 ( .A1(n7303), .A2(n7304), .A3(n7305), .A4(n7306), .ZN(
        vectorData1[50]) );
  AOI22D1BWP U8106 ( .A1(n3576), .A2(\vrf/regTable[5][50] ), .B1(n3595), .B2(
        \vrf/regTable[7][50] ), .ZN(n7306) );
  AOI22D1BWP U8107 ( .A1(n3574), .A2(\vrf/regTable[4][50] ), .B1(n3596), .B2(
        \vrf/regTable[6][50] ), .ZN(n7305) );
  AOI22D1BWP U8108 ( .A1(n3579), .A2(\vrf/regTable[1][50] ), .B1(n3599), .B2(
        \vrf/regTable[3][50] ), .ZN(n7304) );
  AOI22D1BWP U8109 ( .A1(n3581), .A2(\vrf/regTable[0][50] ), .B1(n3594), .B2(
        \vrf/regTable[2][50] ), .ZN(n7303) );
  ND4D1BWP U8110 ( .A1(n8071), .A2(n8072), .A3(n8073), .A4(n8074), .ZN(
        vectorData1[242]) );
  AOI22D1BWP U8111 ( .A1(n3576), .A2(\vrf/regTable[5][242] ), .B1(n3567), .B2(
        \vrf/regTable[7][242] ), .ZN(n8074) );
  AOI22D1BWP U8112 ( .A1(n3574), .A2(\vrf/regTable[4][242] ), .B1(n3570), .B2(
        \vrf/regTable[6][242] ), .ZN(n8073) );
  AOI22D1BWP U8113 ( .A1(n3579), .A2(\vrf/regTable[1][242] ), .B1(n3575), .B2(
        \vrf/regTable[3][242] ), .ZN(n8072) );
  AOI22D1BWP U8114 ( .A1(n3581), .A2(\vrf/regTable[0][242] ), .B1(n3572), .B2(
        \vrf/regTable[2][242] ), .ZN(n8071) );
  AOI22D1BWP U8115 ( .A1(n5231), .A2(vectorData1[114]), .B1(n5184), .B2(
        vectorData1[18]), .ZN(n5025) );
  ND4D1BWP U8116 ( .A1(n7175), .A2(n7176), .A3(n7177), .A4(n7178), .ZN(
        vectorData1[18]) );
  AOI22D1BWP U8117 ( .A1(n3576), .A2(\vrf/regTable[5][18] ), .B1(n3567), .B2(
        \vrf/regTable[7][18] ), .ZN(n7178) );
  AOI22D1BWP U8118 ( .A1(n3574), .A2(\vrf/regTable[4][18] ), .B1(n3570), .B2(
        \vrf/regTable[6][18] ), .ZN(n7177) );
  AOI22D1BWP U8119 ( .A1(n3579), .A2(\vrf/regTable[1][18] ), .B1(n3575), .B2(
        \vrf/regTable[3][18] ), .ZN(n7176) );
  AOI22D1BWP U8120 ( .A1(n3581), .A2(\vrf/regTable[0][18] ), .B1(n3572), .B2(
        \vrf/regTable[2][18] ), .ZN(n7175) );
  ND4D1BWP U8121 ( .A1(n7559), .A2(n7560), .A3(n7561), .A4(n7562), .ZN(
        vectorData1[114]) );
  AOI22D1BWP U8122 ( .A1(n3576), .A2(\vrf/regTable[5][114] ), .B1(n3595), .B2(
        \vrf/regTable[7][114] ), .ZN(n7562) );
  AOI22D1BWP U8123 ( .A1(n3574), .A2(\vrf/regTable[4][114] ), .B1(n3596), .B2(
        \vrf/regTable[6][114] ), .ZN(n7561) );
  AOI22D1BWP U8124 ( .A1(n3579), .A2(\vrf/regTable[1][114] ), .B1(n3599), .B2(
        \vrf/regTable[3][114] ), .ZN(n7560) );
  AOI22D1BWP U8125 ( .A1(n3581), .A2(\vrf/regTable[0][114] ), .B1(n3594), .B2(
        \vrf/regTable[2][114] ), .ZN(n7559) );
  ND4D1BWP U8126 ( .A1(n8297), .A2(n8298), .A3(n8299), .A4(n8300), .ZN(
        scalarData1[2]) );
  AOI22D1BWP U8127 ( .A1(n8287), .A2(\srf/regTable[5][2] ), .B1(n8288), .B2(
        \srf/regTable[7][2] ), .ZN(n8300) );
  AOI22D1BWP U8128 ( .A1(n8285), .A2(\srf/regTable[4][2] ), .B1(n8286), .B2(
        \srf/regTable[6][2] ), .ZN(n8299) );
  AOI22D1BWP U8129 ( .A1(n8282), .A2(\srf/regTable[1][2] ), .B1(n8284), .B2(
        \srf/regTable[3][2] ), .ZN(n8298) );
  AOI22D1BWP U8130 ( .A1(n8278), .A2(\srf/regTable[0][2] ), .B1(n8280), .B2(
        \srf/regTable[2][2] ), .ZN(n8297) );
  OAI211D1BWP U8131 ( .A1(n5497), .A2(n4405), .B(n5359), .C(n4535), .ZN(N4373)
         );
  AOI22D1BWP U8132 ( .A1(n3669), .A2(vectorToLoad[155]), .B1(n4627), .B2(n5358), .ZN(n5359) );
  NR2XD0BWP U8133 ( .A1(n5334), .A2(\intadd_34/A[0] ), .ZN(n5358) );
  NR2XD0BWP U8134 ( .A1(n5278), .A2(cycles[0]), .ZN(n5357) );
  OAI211D1BWP U8135 ( .A1(n5360), .A2(n5509), .B(n5361), .C(n4406), .ZN(N4374)
         );
  AOI22D1BWP U8136 ( .A1(n3668), .A2(vectorToLoad[156]), .B1(n4626), .B2(n5406), .ZN(n5361) );
  NR2XD0BWP U8137 ( .A1(n5279), .A2(cycles[0]), .ZN(n5406) );
  AO222D1BWP U8138 ( .A1(n3642), .A2(n4548), .B1(n5528), .B2(n3667), .C1(n3668), .C2(vectorToLoad[104]), .Z(N4321) );
  NR2XD0BWP U8139 ( .A1(n4652), .A2(n5282), .ZN(n5528) );
  AO211D1BWP U8140 ( .A1(n4073), .A2(scalarData1[1]), .B(n3948), .C(n3947), 
        .Z(N4177) );
  AO22D1BWP U8141 ( .A1(n4072), .A2(vectorData1[1]), .B1(n4071), .B2(Addr[1]), 
        .Z(n3947) );
  ND4D1BWP U8142 ( .A1(n7123), .A2(n7124), .A3(n7125), .A4(n7126), .ZN(
        vectorData1[1]) );
  AOI22D1BWP U8143 ( .A1(n7117), .A2(\vrf/regTable[5][1] ), .B1(n3595), .B2(
        \vrf/regTable[7][1] ), .ZN(n7126) );
  AOI22D1BWP U8144 ( .A1(n3574), .A2(\vrf/regTable[4][1] ), .B1(n3596), .B2(
        \vrf/regTable[6][1] ), .ZN(n7125) );
  AOI22D1BWP U8145 ( .A1(n7112), .A2(\vrf/regTable[1][1] ), .B1(n3599), .B2(
        \vrf/regTable[3][1] ), .ZN(n7124) );
  AOI22D1BWP U8146 ( .A1(n3581), .A2(\vrf/regTable[0][1] ), .B1(n3594), .B2(
        \vrf/regTable[2][1] ), .ZN(n7123) );
  AOI31D1BWP U8147 ( .A1(n5016), .A2(n5015), .A3(n5017), .B(n4070), .ZN(n3948)
         );
  AOI22D1BWP U8148 ( .A1(n5228), .A2(vectorData1[209]), .B1(n5231), .B2(
        vectorData1[113]), .ZN(n5017) );
  ND4D1BWP U8149 ( .A1(n7555), .A2(n7556), .A3(n7557), .A4(n7558), .ZN(
        vectorData1[113]) );
  AOI22D1BWP U8150 ( .A1(n3576), .A2(\vrf/regTable[5][113] ), .B1(n3567), .B2(
        \vrf/regTable[7][113] ), .ZN(n7558) );
  AOI22D1BWP U8151 ( .A1(n3574), .A2(\vrf/regTable[4][113] ), .B1(n3570), .B2(
        \vrf/regTable[6][113] ), .ZN(n7557) );
  AOI22D1BWP U8152 ( .A1(n3579), .A2(\vrf/regTable[1][113] ), .B1(n3599), .B2(
        \vrf/regTable[3][113] ), .ZN(n7556) );
  AOI22D1BWP U8153 ( .A1(n3581), .A2(\vrf/regTable[0][113] ), .B1(n3572), .B2(
        \vrf/regTable[2][113] ), .ZN(n7555) );
  ND4D1BWP U8154 ( .A1(n7939), .A2(n7940), .A3(n7941), .A4(n7942), .ZN(
        vectorData1[209]) );
  AOI22D1BWP U8155 ( .A1(n3576), .A2(\vrf/regTable[5][209] ), .B1(n3567), .B2(
        \vrf/regTable[7][209] ), .ZN(n7942) );
  AOI22D1BWP U8156 ( .A1(n3574), .A2(\vrf/regTable[4][209] ), .B1(n3570), .B2(
        \vrf/regTable[6][209] ), .ZN(n7941) );
  AOI22D1BWP U8157 ( .A1(n3579), .A2(\vrf/regTable[1][209] ), .B1(n3575), .B2(
        \vrf/regTable[3][209] ), .ZN(n7940) );
  AOI22D1BWP U8158 ( .A1(n3581), .A2(\vrf/regTable[0][209] ), .B1(n3572), .B2(
        \vrf/regTable[2][209] ), .ZN(n7939) );
  AOI211XD0BWP U8159 ( .A1(n5185), .A2(vectorData1[81]), .B(n5014), .C(n5013), 
        .ZN(n5015) );
  ND4D1BWP U8160 ( .A1(n5012), .A2(n5011), .A3(n5010), .A4(n5009), .ZN(n5013)
         );
  AOI22D1BWP U8161 ( .A1(n5187), .A2(vectorData1[225]), .B1(n3601), .B2(
        vectorData1[33]), .ZN(n5009) );
  ND4D1BWP U8162 ( .A1(n7235), .A2(n7236), .A3(n7237), .A4(n7238), .ZN(
        vectorData1[33]) );
  AOI22D1BWP U8163 ( .A1(n3576), .A2(\vrf/regTable[5][33] ), .B1(n3567), .B2(
        \vrf/regTable[7][33] ), .ZN(n7238) );
  AOI22D1BWP U8164 ( .A1(n3574), .A2(\vrf/regTable[4][33] ), .B1(n3570), .B2(
        \vrf/regTable[6][33] ), .ZN(n7237) );
  AOI22D1BWP U8165 ( .A1(n3579), .A2(\vrf/regTable[1][33] ), .B1(n3575), .B2(
        \vrf/regTable[3][33] ), .ZN(n7236) );
  AOI22D1BWP U8166 ( .A1(n3581), .A2(\vrf/regTable[0][33] ), .B1(n3572), .B2(
        \vrf/regTable[2][33] ), .ZN(n7235) );
  ND4D1BWP U8167 ( .A1(n8003), .A2(n8004), .A3(n8005), .A4(n8006), .ZN(
        vectorData1[225]) );
  AOI22D1BWP U8168 ( .A1(n3576), .A2(\vrf/regTable[5][225] ), .B1(n3595), .B2(
        \vrf/regTable[7][225] ), .ZN(n8006) );
  AOI22D1BWP U8169 ( .A1(n3574), .A2(\vrf/regTable[4][225] ), .B1(n3596), .B2(
        \vrf/regTable[6][225] ), .ZN(n8005) );
  AOI22D1BWP U8170 ( .A1(n3579), .A2(\vrf/regTable[1][225] ), .B1(n3599), .B2(
        \vrf/regTable[3][225] ), .ZN(n8004) );
  AOI22D1BWP U8171 ( .A1(n3581), .A2(\vrf/regTable[0][225] ), .B1(n3594), .B2(
        \vrf/regTable[2][225] ), .ZN(n8003) );
  AOI22D1BWP U8172 ( .A1(n3671), .A2(vectorData1[97]), .B1(n5186), .B2(
        vectorData1[65]), .ZN(n5010) );
  ND4D1BWP U8173 ( .A1(n7363), .A2(n7364), .A3(n7365), .A4(n7366), .ZN(
        vectorData1[65]) );
  AOI22D1BWP U8174 ( .A1(n3576), .A2(\vrf/regTable[5][65] ), .B1(n3567), .B2(
        \vrf/regTable[7][65] ), .ZN(n7366) );
  AOI22D1BWP U8175 ( .A1(n3574), .A2(\vrf/regTable[4][65] ), .B1(n3570), .B2(
        \vrf/regTable[6][65] ), .ZN(n7365) );
  AOI22D1BWP U8176 ( .A1(n3579), .A2(\vrf/regTable[1][65] ), .B1(n3575), .B2(
        \vrf/regTable[3][65] ), .ZN(n7364) );
  AOI22D1BWP U8177 ( .A1(n3581), .A2(\vrf/regTable[0][65] ), .B1(n3572), .B2(
        \vrf/regTable[2][65] ), .ZN(n7363) );
  ND4D1BWP U8178 ( .A1(n7491), .A2(n7492), .A3(n7493), .A4(n7494), .ZN(
        vectorData1[97]) );
  AOI22D1BWP U8179 ( .A1(n3576), .A2(\vrf/regTable[5][97] ), .B1(n3567), .B2(
        \vrf/regTable[7][97] ), .ZN(n7494) );
  AOI22D1BWP U8180 ( .A1(n3574), .A2(\vrf/regTable[4][97] ), .B1(n3570), .B2(
        \vrf/regTable[6][97] ), .ZN(n7493) );
  AOI22D1BWP U8181 ( .A1(n3579), .A2(\vrf/regTable[1][97] ), .B1(n3575), .B2(
        \vrf/regTable[3][97] ), .ZN(n7492) );
  AOI22D1BWP U8182 ( .A1(n3581), .A2(\vrf/regTable[0][97] ), .B1(n3572), .B2(
        \vrf/regTable[2][97] ), .ZN(n7491) );
  AOI22D1BWP U8183 ( .A1(n5226), .A2(vectorData1[129]), .B1(n5184), .B2(
        vectorData1[17]), .ZN(n5011) );
  ND4D1BWP U8184 ( .A1(n7171), .A2(n7172), .A3(n7173), .A4(n7174), .ZN(
        vectorData1[17]) );
  AOI22D1BWP U8185 ( .A1(n3576), .A2(\vrf/regTable[5][17] ), .B1(n3595), .B2(
        \vrf/regTable[7][17] ), .ZN(n7174) );
  AOI22D1BWP U8186 ( .A1(n3574), .A2(\vrf/regTable[4][17] ), .B1(n3596), .B2(
        \vrf/regTable[6][17] ), .ZN(n7173) );
  AOI22D1BWP U8187 ( .A1(n3579), .A2(\vrf/regTable[1][17] ), .B1(n3599), .B2(
        \vrf/regTable[3][17] ), .ZN(n7172) );
  AOI22D1BWP U8188 ( .A1(n3581), .A2(\vrf/regTable[0][17] ), .B1(n3594), .B2(
        \vrf/regTable[2][17] ), .ZN(n7171) );
  ND4D1BWP U8189 ( .A1(n7619), .A2(n7620), .A3(n7621), .A4(n7622), .ZN(
        vectorData1[129]) );
  AOI22D1BWP U8190 ( .A1(n3576), .A2(\vrf/regTable[5][129] ), .B1(n3567), .B2(
        \vrf/regTable[7][129] ), .ZN(n7622) );
  AOI22D1BWP U8191 ( .A1(n3574), .A2(\vrf/regTable[4][129] ), .B1(n3570), .B2(
        \vrf/regTable[6][129] ), .ZN(n7621) );
  AOI22D1BWP U8192 ( .A1(n3579), .A2(\vrf/regTable[1][129] ), .B1(n3575), .B2(
        \vrf/regTable[3][129] ), .ZN(n7620) );
  AOI22D1BWP U8193 ( .A1(n3581), .A2(\vrf/regTable[0][129] ), .B1(n3572), .B2(
        \vrf/regTable[2][129] ), .ZN(n7619) );
  AOI22D1BWP U8194 ( .A1(n5233), .A2(vectorData1[177]), .B1(n5227), .B2(
        vectorData1[193]), .ZN(n5012) );
  ND4D1BWP U8195 ( .A1(n7875), .A2(n7876), .A3(n7877), .A4(n7878), .ZN(
        vectorData1[193]) );
  AOI22D1BWP U8196 ( .A1(n3576), .A2(\vrf/regTable[5][193] ), .B1(n3595), .B2(
        \vrf/regTable[7][193] ), .ZN(n7878) );
  AOI22D1BWP U8197 ( .A1(n3574), .A2(\vrf/regTable[4][193] ), .B1(n3596), .B2(
        \vrf/regTable[6][193] ), .ZN(n7877) );
  AOI22D1BWP U8198 ( .A1(n3579), .A2(\vrf/regTable[1][193] ), .B1(n3599), .B2(
        \vrf/regTable[3][193] ), .ZN(n7876) );
  AOI22D1BWP U8199 ( .A1(n3581), .A2(\vrf/regTable[0][193] ), .B1(n3594), .B2(
        \vrf/regTable[2][193] ), .ZN(n7875) );
  ND4D1BWP U8200 ( .A1(n7811), .A2(n7812), .A3(n7813), .A4(n7814), .ZN(
        vectorData1[177]) );
  AOI22D1BWP U8201 ( .A1(n3576), .A2(\vrf/regTable[5][177] ), .B1(n3567), .B2(
        \vrf/regTable[7][177] ), .ZN(n7814) );
  AOI22D1BWP U8202 ( .A1(n3574), .A2(\vrf/regTable[4][177] ), .B1(n3570), .B2(
        \vrf/regTable[6][177] ), .ZN(n7813) );
  AOI22D1BWP U8203 ( .A1(n3579), .A2(\vrf/regTable[1][177] ), .B1(n3575), .B2(
        \vrf/regTable[3][177] ), .ZN(n7812) );
  AOI22D1BWP U8204 ( .A1(n3581), .A2(\vrf/regTable[0][177] ), .B1(n3572), .B2(
        \vrf/regTable[2][177] ), .ZN(n7811) );
  AO22D1BWP U8205 ( .A1(n5188), .A2(vectorData1[49]), .B1(n5232), .B2(
        vectorData1[145]), .Z(n5014) );
  ND4D1BWP U8206 ( .A1(n7683), .A2(n7684), .A3(n7685), .A4(n7686), .ZN(
        vectorData1[145]) );
  AOI22D1BWP U8207 ( .A1(n3576), .A2(\vrf/regTable[5][145] ), .B1(n3595), .B2(
        \vrf/regTable[7][145] ), .ZN(n7686) );
  AOI22D1BWP U8208 ( .A1(n3574), .A2(\vrf/regTable[4][145] ), .B1(n3596), .B2(
        \vrf/regTable[6][145] ), .ZN(n7685) );
  AOI22D1BWP U8209 ( .A1(n3579), .A2(\vrf/regTable[1][145] ), .B1(n3599), .B2(
        \vrf/regTable[3][145] ), .ZN(n7684) );
  AOI22D1BWP U8210 ( .A1(n3581), .A2(\vrf/regTable[0][145] ), .B1(n3594), .B2(
        \vrf/regTable[2][145] ), .ZN(n7683) );
  ND4D1BWP U8211 ( .A1(n7299), .A2(n7300), .A3(n7301), .A4(n7302), .ZN(
        vectorData1[49]) );
  AOI22D1BWP U8212 ( .A1(n3576), .A2(\vrf/regTable[5][49] ), .B1(n3595), .B2(
        \vrf/regTable[7][49] ), .ZN(n7302) );
  AOI22D1BWP U8213 ( .A1(n3574), .A2(\vrf/regTable[4][49] ), .B1(n3596), .B2(
        \vrf/regTable[6][49] ), .ZN(n7301) );
  AOI22D1BWP U8214 ( .A1(n3579), .A2(\vrf/regTable[1][49] ), .B1(n3599), .B2(
        \vrf/regTable[3][49] ), .ZN(n7300) );
  AOI22D1BWP U8215 ( .A1(n3581), .A2(\vrf/regTable[0][49] ), .B1(n3594), .B2(
        \vrf/regTable[2][49] ), .ZN(n7299) );
  ND4D1BWP U8216 ( .A1(n7427), .A2(n7428), .A3(n7429), .A4(n7430), .ZN(
        vectorData1[81]) );
  AOI22D1BWP U8217 ( .A1(n3576), .A2(\vrf/regTable[5][81] ), .B1(n3567), .B2(
        \vrf/regTable[7][81] ), .ZN(n7430) );
  AOI22D1BWP U8218 ( .A1(n3574), .A2(\vrf/regTable[4][81] ), .B1(n3570), .B2(
        \vrf/regTable[6][81] ), .ZN(n7429) );
  AOI22D1BWP U8219 ( .A1(n3579), .A2(\vrf/regTable[1][81] ), .B1(n3575), .B2(
        \vrf/regTable[3][81] ), .ZN(n7428) );
  AOI22D1BWP U8220 ( .A1(n3581), .A2(\vrf/regTable[0][81] ), .B1(n3572), .B2(
        \vrf/regTable[2][81] ), .ZN(n7427) );
  AOI22D1BWP U8221 ( .A1(n5229), .A2(vectorData1[241]), .B1(n5230), .B2(
        vectorData1[161]), .ZN(n5016) );
  ND4D1BWP U8222 ( .A1(n7747), .A2(n7748), .A3(n7749), .A4(n7750), .ZN(
        vectorData1[161]) );
  AOI22D1BWP U8223 ( .A1(n3576), .A2(\vrf/regTable[5][161] ), .B1(n3567), .B2(
        \vrf/regTable[7][161] ), .ZN(n7750) );
  AOI22D1BWP U8224 ( .A1(n3574), .A2(\vrf/regTable[4][161] ), .B1(n3570), .B2(
        \vrf/regTable[6][161] ), .ZN(n7749) );
  AOI22D1BWP U8225 ( .A1(n3579), .A2(\vrf/regTable[1][161] ), .B1(n3575), .B2(
        \vrf/regTable[3][161] ), .ZN(n7748) );
  AOI22D1BWP U8226 ( .A1(n3581), .A2(\vrf/regTable[0][161] ), .B1(n3572), .B2(
        \vrf/regTable[2][161] ), .ZN(n7747) );
  ND4D1BWP U8227 ( .A1(n8067), .A2(n8068), .A3(n8069), .A4(n8070), .ZN(
        vectorData1[241]) );
  AOI22D1BWP U8228 ( .A1(n3576), .A2(\vrf/regTable[5][241] ), .B1(n3567), .B2(
        \vrf/regTable[7][241] ), .ZN(n8070) );
  AOI22D1BWP U8229 ( .A1(n3574), .A2(\vrf/regTable[4][241] ), .B1(n3570), .B2(
        \vrf/regTable[6][241] ), .ZN(n8069) );
  AOI22D1BWP U8230 ( .A1(n3579), .A2(\vrf/regTable[1][241] ), .B1(n3575), .B2(
        \vrf/regTable[3][241] ), .ZN(n8068) );
  AOI22D1BWP U8231 ( .A1(n3581), .A2(\vrf/regTable[0][241] ), .B1(n3572), .B2(
        \vrf/regTable[2][241] ), .ZN(n8067) );
  ND4D1BWP U8232 ( .A1(n8293), .A2(n8294), .A3(n8295), .A4(n8296), .ZN(
        scalarData1[1]) );
  AOI22D1BWP U8233 ( .A1(n8287), .A2(\srf/regTable[5][1] ), .B1(n8288), .B2(
        \srf/regTable[7][1] ), .ZN(n8296) );
  AOI22D1BWP U8234 ( .A1(n8285), .A2(\srf/regTable[4][1] ), .B1(n8286), .B2(
        \srf/regTable[6][1] ), .ZN(n8295) );
  AOI22D1BWP U8235 ( .A1(n8282), .A2(\srf/regTable[1][1] ), .B1(n8284), .B2(
        \srf/regTable[3][1] ), .ZN(n8294) );
  AOI22D1BWP U8236 ( .A1(n8278), .A2(\srf/regTable[0][1] ), .B1(n8280), .B2(
        \srf/regTable[2][1] ), .ZN(n8293) );
  OAI211D1BWP U8237 ( .A1(n5362), .A2(n5509), .B(n5363), .C(n4406), .ZN(N4375)
         );
  AOI22D1BWP U8238 ( .A1(n3669), .A2(vectorToLoad[157]), .B1(n4626), .B2(n5408), .ZN(n5363) );
  AO222D1BWP U8239 ( .A1(n3668), .A2(vectorToLoad[47]), .B1(n4549), .B2(n5535), 
        .C1(n3649), .C2(n5330), .Z(N4264) );
  NR2XD0BWP U8240 ( .A1(n3679), .A2(n5283), .ZN(n5330) );
  NR2XD0BWP U8241 ( .A1(n6037), .A2(n5282), .ZN(n5535) );
  OAI211D1BWP U8242 ( .A1(n5364), .A2(n5509), .B(n5365), .C(n4406), .ZN(N4376)
         );
  AOI22D1BWP U8243 ( .A1(n3668), .A2(vectorToLoad[158]), .B1(n4626), .B2(n5410), .ZN(n5365) );
  NR2XD0BWP U8244 ( .A1(n5281), .A2(cycles[0]), .ZN(n5410) );
  AO211D1BWP U8245 ( .A1(n4073), .A2(scalarData1[0]), .B(n3791), .C(n3790), 
        .Z(N4176) );
  MOAI22D0BWP U8246 ( .A1(n3830), .A2(n3789), .B1(n4072), .B2(vectorData1[0]), 
        .ZN(n3790) );
  ND4D1BWP U8247 ( .A1(n7119), .A2(n7120), .A3(n7121), .A4(n7122), .ZN(
        vectorData1[0]) );
  AOI22D1BWP U8248 ( .A1(n3576), .A2(\vrf/regTable[5][0] ), .B1(n3595), .B2(
        \vrf/regTable[7][0] ), .ZN(n7122) );
  AOI22D1BWP U8249 ( .A1(n3574), .A2(\vrf/regTable[4][0] ), .B1(n3596), .B2(
        \vrf/regTable[6][0] ), .ZN(n7121) );
  AOI22D1BWP U8250 ( .A1(n3579), .A2(\vrf/regTable[1][0] ), .B1(n3599), .B2(
        \vrf/regTable[3][0] ), .ZN(n7120) );
  AOI22D1BWP U8251 ( .A1(n3581), .A2(\vrf/regTable[0][0] ), .B1(n3594), .B2(
        \vrf/regTable[2][0] ), .ZN(n7119) );
  AOI31D1BWP U8252 ( .A1(n5007), .A2(n5006), .A3(n5008), .B(n4070), .ZN(n3791)
         );
  AOI22D1BWP U8253 ( .A1(n5231), .A2(vectorData1[112]), .B1(n5185), .B2(
        vectorData1[80]), .ZN(n5008) );
  ND4D1BWP U8254 ( .A1(n7423), .A2(n7424), .A3(n7425), .A4(n7426), .ZN(
        vectorData1[80]) );
  AOI22D1BWP U8255 ( .A1(n3576), .A2(\vrf/regTable[5][80] ), .B1(n3567), .B2(
        \vrf/regTable[7][80] ), .ZN(n7426) );
  AOI22D1BWP U8256 ( .A1(n3574), .A2(\vrf/regTable[4][80] ), .B1(n3570), .B2(
        \vrf/regTable[6][80] ), .ZN(n7425) );
  AOI22D1BWP U8257 ( .A1(n3579), .A2(\vrf/regTable[1][80] ), .B1(n3575), .B2(
        \vrf/regTable[3][80] ), .ZN(n7424) );
  AOI22D1BWP U8258 ( .A1(n3581), .A2(\vrf/regTable[0][80] ), .B1(n3572), .B2(
        \vrf/regTable[2][80] ), .ZN(n7423) );
  ND4D1BWP U8259 ( .A1(n7551), .A2(n7552), .A3(n7553), .A4(n7554), .ZN(
        vectorData1[112]) );
  AOI22D1BWP U8260 ( .A1(n3576), .A2(\vrf/regTable[5][112] ), .B1(n3595), .B2(
        \vrf/regTable[7][112] ), .ZN(n7554) );
  AOI22D1BWP U8261 ( .A1(n3574), .A2(\vrf/regTable[4][112] ), .B1(n3596), .B2(
        \vrf/regTable[6][112] ), .ZN(n7553) );
  AOI22D1BWP U8262 ( .A1(n3579), .A2(\vrf/regTable[1][112] ), .B1(n3599), .B2(
        \vrf/regTable[3][112] ), .ZN(n7552) );
  AOI22D1BWP U8263 ( .A1(n3581), .A2(\vrf/regTable[0][112] ), .B1(n3594), .B2(
        \vrf/regTable[2][112] ), .ZN(n7551) );
  AOI211XD0BWP U8264 ( .A1(n5226), .A2(vectorData1[128]), .B(n5005), .C(n5004), 
        .ZN(n5006) );
  ND4D1BWP U8265 ( .A1(n5003), .A2(n5002), .A3(n5001), .A4(n5000), .ZN(n5004)
         );
  AOI22D1BWP U8266 ( .A1(n5232), .A2(vectorData1[144]), .B1(n5230), .B2(
        vectorData1[160]), .ZN(n5000) );
  ND4D1BWP U8267 ( .A1(n7743), .A2(n7744), .A3(n7745), .A4(n7746), .ZN(
        vectorData1[160]) );
  AOI22D1BWP U8268 ( .A1(n3576), .A2(\vrf/regTable[5][160] ), .B1(n3595), .B2(
        \vrf/regTable[7][160] ), .ZN(n7746) );
  AOI22D1BWP U8269 ( .A1(n3574), .A2(\vrf/regTable[4][160] ), .B1(n3596), .B2(
        \vrf/regTable[6][160] ), .ZN(n7745) );
  AOI22D1BWP U8270 ( .A1(n3579), .A2(\vrf/regTable[1][160] ), .B1(n3575), .B2(
        \vrf/regTable[3][160] ), .ZN(n7744) );
  AOI22D1BWP U8271 ( .A1(n3581), .A2(\vrf/regTable[0][160] ), .B1(n3594), .B2(
        \vrf/regTable[2][160] ), .ZN(n7743) );
  ND4D1BWP U8272 ( .A1(n7679), .A2(n7680), .A3(n7681), .A4(n7682), .ZN(
        vectorData1[144]) );
  AOI22D1BWP U8273 ( .A1(n3576), .A2(\vrf/regTable[5][144] ), .B1(n3595), .B2(
        \vrf/regTable[7][144] ), .ZN(n7682) );
  AOI22D1BWP U8274 ( .A1(n3574), .A2(\vrf/regTable[4][144] ), .B1(n3596), .B2(
        \vrf/regTable[6][144] ), .ZN(n7681) );
  AOI22D1BWP U8275 ( .A1(n3579), .A2(\vrf/regTable[1][144] ), .B1(n3599), .B2(
        \vrf/regTable[3][144] ), .ZN(n7680) );
  AOI22D1BWP U8276 ( .A1(n3581), .A2(\vrf/regTable[0][144] ), .B1(n3594), .B2(
        \vrf/regTable[2][144] ), .ZN(n7679) );
  AOI22D1BWP U8277 ( .A1(n5186), .A2(vectorData1[64]), .B1(n5227), .B2(
        vectorData1[192]), .ZN(n5001) );
  ND4D1BWP U8278 ( .A1(n7871), .A2(n7872), .A3(n7873), .A4(n7874), .ZN(
        vectorData1[192]) );
  AOI22D1BWP U8279 ( .A1(n3576), .A2(\vrf/regTable[5][192] ), .B1(n3595), .B2(
        \vrf/regTable[7][192] ), .ZN(n7874) );
  AOI22D1BWP U8280 ( .A1(n3574), .A2(\vrf/regTable[4][192] ), .B1(n3596), .B2(
        \vrf/regTable[6][192] ), .ZN(n7873) );
  AOI22D1BWP U8281 ( .A1(n3579), .A2(\vrf/regTable[1][192] ), .B1(n3599), .B2(
        \vrf/regTable[3][192] ), .ZN(n7872) );
  AOI22D1BWP U8282 ( .A1(n3581), .A2(\vrf/regTable[0][192] ), .B1(n3594), .B2(
        \vrf/regTable[2][192] ), .ZN(n7871) );
  ND4D1BWP U8283 ( .A1(n7359), .A2(n7360), .A3(n7361), .A4(n7362), .ZN(
        vectorData1[64]) );
  AOI22D1BWP U8284 ( .A1(n3576), .A2(\vrf/regTable[5][64] ), .B1(n3595), .B2(
        \vrf/regTable[7][64] ), .ZN(n7362) );
  AOI22D1BWP U8285 ( .A1(n3574), .A2(\vrf/regTable[4][64] ), .B1(n3596), .B2(
        \vrf/regTable[6][64] ), .ZN(n7361) );
  AOI22D1BWP U8286 ( .A1(n3579), .A2(\vrf/regTable[1][64] ), .B1(n3599), .B2(
        \vrf/regTable[3][64] ), .ZN(n7360) );
  AOI22D1BWP U8287 ( .A1(n3581), .A2(\vrf/regTable[0][64] ), .B1(n3594), .B2(
        \vrf/regTable[2][64] ), .ZN(n7359) );
  AOI22D1BWP U8288 ( .A1(n5233), .A2(vectorData1[176]), .B1(n3601), .B2(
        vectorData1[32]), .ZN(n5002) );
  ND4D1BWP U8289 ( .A1(n7231), .A2(n7232), .A3(n7233), .A4(n7234), .ZN(
        vectorData1[32]) );
  AOI22D1BWP U8290 ( .A1(n3576), .A2(\vrf/regTable[5][32] ), .B1(n3595), .B2(
        \vrf/regTable[7][32] ), .ZN(n7234) );
  AOI22D1BWP U8291 ( .A1(n3574), .A2(\vrf/regTable[4][32] ), .B1(n3596), .B2(
        \vrf/regTable[6][32] ), .ZN(n7233) );
  AOI22D1BWP U8292 ( .A1(n3579), .A2(\vrf/regTable[1][32] ), .B1(n3599), .B2(
        \vrf/regTable[3][32] ), .ZN(n7232) );
  AOI22D1BWP U8293 ( .A1(n3581), .A2(\vrf/regTable[0][32] ), .B1(n3594), .B2(
        \vrf/regTable[2][32] ), .ZN(n7231) );
  ND4D1BWP U8294 ( .A1(n7807), .A2(n7808), .A3(n7809), .A4(n7810), .ZN(
        vectorData1[176]) );
  AOI22D1BWP U8295 ( .A1(n3576), .A2(\vrf/regTable[5][176] ), .B1(n3595), .B2(
        \vrf/regTable[7][176] ), .ZN(n7810) );
  AOI22D1BWP U8296 ( .A1(n3574), .A2(\vrf/regTable[4][176] ), .B1(n3596), .B2(
        \vrf/regTable[6][176] ), .ZN(n7809) );
  AOI22D1BWP U8297 ( .A1(n3579), .A2(\vrf/regTable[1][176] ), .B1(n3599), .B2(
        \vrf/regTable[3][176] ), .ZN(n7808) );
  AOI22D1BWP U8298 ( .A1(n3581), .A2(\vrf/regTable[0][176] ), .B1(n3594), .B2(
        \vrf/regTable[2][176] ), .ZN(n7807) );
  AOI22D1BWP U8299 ( .A1(n5188), .A2(vectorData1[48]), .B1(n5184), .B2(
        vectorData1[16]), .ZN(n5003) );
  ND4D1BWP U8300 ( .A1(n7167), .A2(n7168), .A3(n7169), .A4(n7170), .ZN(
        vectorData1[16]) );
  AOI22D1BWP U8301 ( .A1(n3576), .A2(\vrf/regTable[5][16] ), .B1(n3567), .B2(
        \vrf/regTable[7][16] ), .ZN(n7170) );
  AOI22D1BWP U8302 ( .A1(n3574), .A2(\vrf/regTable[4][16] ), .B1(n3570), .B2(
        \vrf/regTable[6][16] ), .ZN(n7169) );
  AOI22D1BWP U8303 ( .A1(n3579), .A2(\vrf/regTable[1][16] ), .B1(n3575), .B2(
        \vrf/regTable[3][16] ), .ZN(n7168) );
  AOI22D1BWP U8304 ( .A1(n3581), .A2(\vrf/regTable[0][16] ), .B1(n3572), .B2(
        \vrf/regTable[2][16] ), .ZN(n7167) );
  ND4D1BWP U8305 ( .A1(n7295), .A2(n7296), .A3(n7297), .A4(n7298), .ZN(
        vectorData1[48]) );
  AOI22D1BWP U8306 ( .A1(n3576), .A2(\vrf/regTable[5][48] ), .B1(n3595), .B2(
        \vrf/regTable[7][48] ), .ZN(n7298) );
  AOI22D1BWP U8307 ( .A1(n3574), .A2(\vrf/regTable[4][48] ), .B1(n3596), .B2(
        \vrf/regTable[6][48] ), .ZN(n7297) );
  AOI22D1BWP U8308 ( .A1(n3579), .A2(\vrf/regTable[1][48] ), .B1(n3599), .B2(
        \vrf/regTable[3][48] ), .ZN(n7296) );
  AOI22D1BWP U8309 ( .A1(n3581), .A2(\vrf/regTable[0][48] ), .B1(n3594), .B2(
        \vrf/regTable[2][48] ), .ZN(n7295) );
  AO22D1BWP U8310 ( .A1(n3671), .A2(vectorData1[96]), .B1(n5229), .B2(
        vectorData1[240]), .Z(n5005) );
  ND4D1BWP U8311 ( .A1(n8063), .A2(n8064), .A3(n8065), .A4(n8066), .ZN(
        vectorData1[240]) );
  AOI22D1BWP U8312 ( .A1(n3576), .A2(\vrf/regTable[5][240] ), .B1(n3567), .B2(
        \vrf/regTable[7][240] ), .ZN(n8066) );
  AOI22D1BWP U8313 ( .A1(n3574), .A2(\vrf/regTable[4][240] ), .B1(n3570), .B2(
        \vrf/regTable[6][240] ), .ZN(n8065) );
  AOI22D1BWP U8314 ( .A1(n3579), .A2(\vrf/regTable[1][240] ), .B1(n3575), .B2(
        \vrf/regTable[3][240] ), .ZN(n8064) );
  AOI22D1BWP U8315 ( .A1(n3581), .A2(\vrf/regTable[0][240] ), .B1(n3572), .B2(
        \vrf/regTable[2][240] ), .ZN(n8063) );
  ND4D1BWP U8316 ( .A1(n7487), .A2(n7488), .A3(n7489), .A4(n7490), .ZN(
        vectorData1[96]) );
  AOI22D1BWP U8317 ( .A1(n3576), .A2(\vrf/regTable[5][96] ), .B1(n3567), .B2(
        \vrf/regTable[7][96] ), .ZN(n7490) );
  AOI22D1BWP U8318 ( .A1(n7115), .A2(\vrf/regTable[4][96] ), .B1(n3570), .B2(
        \vrf/regTable[6][96] ), .ZN(n7489) );
  AOI22D1BWP U8319 ( .A1(n3579), .A2(\vrf/regTable[1][96] ), .B1(n3575), .B2(
        \vrf/regTable[3][96] ), .ZN(n7488) );
  AOI22D1BWP U8320 ( .A1(n7108), .A2(\vrf/regTable[0][96] ), .B1(n3572), .B2(
        \vrf/regTable[2][96] ), .ZN(n7487) );
  ND4D1BWP U8321 ( .A1(n7615), .A2(n7616), .A3(n7617), .A4(n7618), .ZN(
        vectorData1[128]) );
  AOI22D1BWP U8322 ( .A1(n3576), .A2(\vrf/regTable[5][128] ), .B1(n3567), .B2(
        \vrf/regTable[7][128] ), .ZN(n7618) );
  AOI22D1BWP U8323 ( .A1(n3574), .A2(\vrf/regTable[4][128] ), .B1(n3570), .B2(
        \vrf/regTable[6][128] ), .ZN(n7617) );
  AOI22D1BWP U8324 ( .A1(n3579), .A2(\vrf/regTable[1][128] ), .B1(n3599), .B2(
        \vrf/regTable[3][128] ), .ZN(n7616) );
  AOI22D1BWP U8325 ( .A1(n3581), .A2(\vrf/regTable[0][128] ), .B1(n3572), .B2(
        \vrf/regTable[2][128] ), .ZN(n7615) );
  AOI22D1BWP U8326 ( .A1(n5228), .A2(vectorData1[208]), .B1(n5187), .B2(
        vectorData1[224]), .ZN(n5007) );
  ND4D1BWP U8327 ( .A1(n7999), .A2(n8000), .A3(n8001), .A4(n8002), .ZN(
        vectorData1[224]) );
  AOI22D1BWP U8328 ( .A1(n3576), .A2(\vrf/regTable[5][224] ), .B1(n3567), .B2(
        \vrf/regTable[7][224] ), .ZN(n8002) );
  AOI22D1BWP U8329 ( .A1(n3574), .A2(\vrf/regTable[4][224] ), .B1(n3570), .B2(
        \vrf/regTable[6][224] ), .ZN(n8001) );
  AOI22D1BWP U8330 ( .A1(n3579), .A2(\vrf/regTable[1][224] ), .B1(n3575), .B2(
        \vrf/regTable[3][224] ), .ZN(n8000) );
  AOI22D1BWP U8331 ( .A1(n3581), .A2(\vrf/regTable[0][224] ), .B1(n3572), .B2(
        \vrf/regTable[2][224] ), .ZN(n7999) );
  ND4D1BWP U8332 ( .A1(n7935), .A2(n7936), .A3(n7937), .A4(n7938), .ZN(
        vectorData1[208]) );
  AOI22D1BWP U8333 ( .A1(n3576), .A2(\vrf/regTable[5][208] ), .B1(n3567), .B2(
        \vrf/regTable[7][208] ), .ZN(n7938) );
  AOI22D1BWP U8334 ( .A1(n3574), .A2(\vrf/regTable[4][208] ), .B1(n3570), .B2(
        \vrf/regTable[6][208] ), .ZN(n7937) );
  AOI22D1BWP U8335 ( .A1(n3579), .A2(\vrf/regTable[1][208] ), .B1(n3575), .B2(
        \vrf/regTable[3][208] ), .ZN(n7936) );
  AOI22D1BWP U8336 ( .A1(n3581), .A2(\vrf/regTable[0][208] ), .B1(n3572), .B2(
        \vrf/regTable[2][208] ), .ZN(n7935) );
  ND4D1BWP U8337 ( .A1(n8289), .A2(n8290), .A3(n8291), .A4(n8292), .ZN(
        scalarData1[0]) );
  AOI22D1BWP U8338 ( .A1(n8287), .A2(\srf/regTable[5][0] ), .B1(n8288), .B2(
        \srf/regTable[7][0] ), .ZN(n8292) );
  AOI22D1BWP U8339 ( .A1(n8285), .A2(\srf/regTable[4][0] ), .B1(n8286), .B2(
        \srf/regTable[6][0] ), .ZN(n8291) );
  AOI22D1BWP U8340 ( .A1(n8282), .A2(\srf/regTable[1][0] ), .B1(n8284), .B2(
        \srf/regTable[3][0] ), .ZN(n8290) );
  AOI22D1BWP U8341 ( .A1(n8278), .A2(\srf/regTable[0][0] ), .B1(n8280), .B2(
        \srf/regTable[2][0] ), .ZN(n8289) );
  OAI211D1BWP U8342 ( .A1(n5366), .A2(n5509), .B(n5367), .C(n4406), .ZN(N4377)
         );
  AOI22D1BWP U8343 ( .A1(n3669), .A2(vectorToLoad[159]), .B1(n4626), .B2(n5412), .ZN(n5367) );
  NR2XD0BWP U8344 ( .A1(n5283), .A2(cycles[0]), .ZN(n5412) );
  OAI211D1BWP U8345 ( .A1(n5370), .A2(n4407), .B(n5369), .C(n4535), .ZN(N4378)
         );
  AOI22D1BWP U8346 ( .A1(n3668), .A2(vectorToLoad[160]), .B1(n5415), .B2(n5511), .ZN(n5369) );
  OAI32D1BWP U8347 ( .A1(n5267), .A2(n5286), .A3(n3679), .B1(n136), .B2(n5267), 
        .ZN(n5511) );
  NR2XD0BWP U8348 ( .A1(n5417), .A2(n5418), .ZN(n5267) );
  AO31D1BWP U8349 ( .A1(n156), .A2(overflow), .A3(n4572), .B(n5247), .Z(N4210)
         );
  AO222D1BWP U8350 ( .A1(n3669), .A2(vectorToLoad[46]), .B1(n4549), .B2(n5534), 
        .C1(n3649), .C2(n5328), .Z(N4263) );
  NR2XD0BWP U8351 ( .A1(\intadd_34/A[3] ), .A2(n5282), .ZN(n5534) );
  OAI211D1BWP U8352 ( .A1(n5517), .A2(n4407), .B(n5371), .C(n4535), .ZN(N4379)
         );
  AOI22D1BWP U8353 ( .A1(n3669), .A2(vectorToLoad[161]), .B1(n5415), .B2(n5515), .ZN(n5371) );
  NR2XD0BWP U8354 ( .A1(n4643), .A2(n5282), .ZN(n5515) );
  OAI211D1BWP U8355 ( .A1(n5520), .A2(n4407), .B(n5372), .C(n4535), .ZN(N4380)
         );
  AOI22D1BWP U8356 ( .A1(n3668), .A2(vectorToLoad[162]), .B1(n5415), .B2(n5518), .ZN(n5372) );
  NR2XD0BWP U8357 ( .A1(n4668), .A2(n5282), .ZN(n5518) );
  AO222D1BWP U8358 ( .A1(n3643), .A2(n4548), .B1(n5529), .B2(n3667), .C1(n3668), .C2(vectorToLoad[105]), .Z(N4322) );
  NR2XD0BWP U8359 ( .A1(n4651), .A2(n5282), .ZN(n5529) );
  OAI211D1BWP U8360 ( .A1(n5523), .A2(n4407), .B(n5373), .C(n4535), .ZN(N4381)
         );
  AOI22D1BWP U8361 ( .A1(n3669), .A2(vectorToLoad[163]), .B1(n5415), .B2(n5521), .ZN(n5373) );
  NR2XD0BWP U8362 ( .A1(n6011), .A2(n5282), .ZN(n5521) );
  AO222D1BWP U8363 ( .A1(n3669), .A2(vectorToLoad[45]), .B1(n4549), .B2(n5533), 
        .C1(n3649), .C2(n5326), .Z(N4262) );
  NR2XD0BWP U8364 ( .A1(n3679), .A2(n5280), .ZN(n5326) );
  NR2XD0BWP U8365 ( .A1(\intadd_34/A[2] ), .A2(n5282), .ZN(n5533) );
  OAI211D1BWP U8366 ( .A1(n5428), .A2(n4407), .B(n5374), .C(n4535), .ZN(N4382)
         );
  AOI22D1BWP U8367 ( .A1(n3668), .A2(vectorToLoad[164]), .B1(n5415), .B2(n5524), .ZN(n5374) );
  NR2XD0BWP U8368 ( .A1(n4665), .A2(n5282), .ZN(n5524) );
  OAI211D1BWP U8369 ( .A1(n5431), .A2(n4407), .B(n5375), .C(n4535), .ZN(N4383)
         );
  AOI22D1BWP U8370 ( .A1(n3669), .A2(vectorToLoad[165]), .B1(n5415), .B2(n5525), .ZN(n5375) );
  NR2XD0BWP U8371 ( .A1(n4664), .A2(n5282), .ZN(n5525) );
  OAI211D1BWP U8372 ( .A1(n5503), .A2(n4407), .B(n5409), .C(n4535), .ZN(N4407)
         );
  AOI22D1BWP U8373 ( .A1(n3668), .A2(vectorToLoad[189]), .B1(n5415), .B2(n5551), .ZN(n5409) );
  NR2XD0BWP U8374 ( .A1(n5280), .A2(cycles[0]), .ZN(n5408) );
  OAI22D1BWP U8375 ( .A1(n4967), .A2(n4926), .B1(n4925), .B2(n4962), .ZN(N1822) );
  AOI211XD0BWP U8376 ( .A1(n4956), .A2(n4934), .B(n4924), .C(n4923), .ZN(n4925) );
  OA211D1BWP U8377 ( .A1(n4934), .A2(n4922), .B(n4955), .C(n4964), .Z(n4923)
         );
  NR2XD0BWP U8378 ( .A1(n5249), .A2(result[12]), .ZN(n4926) );
  AOI211XD0BWP U8379 ( .A1(n3944), .A2(instrIn[8]), .B(n3909), .C(n5200), .ZN(
        n3910) );
  AOI31D1BWP U8380 ( .A1(n5173), .A2(n5172), .A3(n5174), .B(n3661), .ZN(n3909)
         );
  AOI22D1BWP U8381 ( .A1(vectorData2[200]), .A2(n5227), .B1(vectorData2[88]), 
        .B2(n5185), .ZN(n5174) );
  AOI211XD0BWP U8382 ( .A1(vectorData2[136]), .A2(n5226), .B(n5171), .C(n5170), 
        .ZN(n5172) );
  ND4D1BWP U8383 ( .A1(n5169), .A2(n5168), .A3(n5167), .A4(n5166), .ZN(n5170)
         );
  AOI22D1BWP U8384 ( .A1(vectorData2[72]), .A2(n5186), .B1(vectorData2[40]), 
        .B2(n3601), .ZN(n5166) );
  AOI22D1BWP U8385 ( .A1(vectorData2[24]), .A2(n5184), .B1(vectorData2[56]), 
        .B2(n5188), .ZN(n5167) );
  AOI22D1BWP U8386 ( .A1(vectorData2[104]), .A2(n3671), .B1(vectorData2[184]), 
        .B2(n5233), .ZN(n5168) );
  AOI22D1BWP U8387 ( .A1(vectorData2[168]), .A2(n5230), .B1(vectorData2[232]), 
        .B2(n5187), .ZN(n5169) );
  AO22D1BWP U8388 ( .A1(vectorData2[216]), .A2(n5228), .B1(vectorData2[248]), 
        .B2(n5229), .Z(n5171) );
  AOI22D1BWP U8389 ( .A1(vectorData2[152]), .A2(n5232), .B1(vectorData2[120]), 
        .B2(n5231), .ZN(n5173) );
  AOI22D1BWP U8390 ( .A1(n4681), .A2(vectorData2[8]), .B1(n4688), .B2(
        scalarData2[8]), .ZN(n3911) );
  OAI211D1BWP U8391 ( .A1(n3844), .A2(n153), .B(n3843), .C(n3842), .ZN(N4197)
         );
  AOI21D1BWP U8392 ( .A1(scalarData2[5]), .A2(n4688), .B(n3841), .ZN(n3843) );
  AOI31D1BWP U8393 ( .A1(n5164), .A2(n5163), .A3(n5165), .B(n3661), .ZN(n3841)
         );
  AOI22D1BWP U8394 ( .A1(vectorData2[213]), .A2(n5228), .B1(vectorData2[197]), 
        .B2(n5227), .ZN(n5165) );
  AOI211XD0BWP U8395 ( .A1(vectorData2[149]), .A2(n5232), .B(n5162), .C(n5161), 
        .ZN(n5163) );
  ND4D1BWP U8396 ( .A1(n5160), .A2(n5159), .A3(n5158), .A4(n5157), .ZN(n5161)
         );
  AOI22D1BWP U8397 ( .A1(vectorData2[53]), .A2(n5188), .B1(vectorData2[117]), 
        .B2(n5231), .ZN(n5157) );
  AOI22D1BWP U8398 ( .A1(vectorData2[37]), .A2(n3601), .B1(vectorData2[165]), 
        .B2(n5230), .ZN(n5158) );
  AOI22D1BWP U8399 ( .A1(vectorData2[133]), .A2(n5226), .B1(vectorData2[229]), 
        .B2(n5187), .ZN(n5159) );
  AOI22D1BWP U8400 ( .A1(vectorData2[101]), .A2(n3671), .B1(vectorData2[69]), 
        .B2(n5186), .ZN(n5160) );
  AO22D1BWP U8401 ( .A1(vectorData2[85]), .A2(n5185), .B1(vectorData2[181]), 
        .B2(n5233), .Z(n5162) );
  AOI22D1BWP U8402 ( .A1(vectorData2[245]), .A2(n5229), .B1(vectorData2[21]), 
        .B2(n5184), .ZN(n5164) );
  AOI211XD0BWP U8403 ( .A1(n3944), .A2(instrIn[9]), .B(n3943), .C(n5200), .ZN(
        n3945) );
  AOI31D1BWP U8404 ( .A1(n5182), .A2(n5181), .A3(n5183), .B(n3661), .ZN(n3943)
         );
  AOI22D1BWP U8405 ( .A1(vectorData2[169]), .A2(n5230), .B1(vectorData2[121]), 
        .B2(n5231), .ZN(n5183) );
  AOI211XD0BWP U8406 ( .A1(vectorData2[57]), .A2(n5188), .B(n5180), .C(n5179), 
        .ZN(n5181) );
  ND4D1BWP U8407 ( .A1(n5178), .A2(n5177), .A3(n5176), .A4(n5175), .ZN(n5179)
         );
  AOI22D1BWP U8408 ( .A1(vectorData2[89]), .A2(n5185), .B1(vectorData2[25]), 
        .B2(n5184), .ZN(n5175) );
  AOI22D1BWP U8409 ( .A1(vectorData2[201]), .A2(n5227), .B1(vectorData2[217]), 
        .B2(n5228), .ZN(n5176) );
  AOI22D1BWP U8410 ( .A1(vectorData2[105]), .A2(n3671), .B1(vectorData2[233]), 
        .B2(n5187), .ZN(n5177) );
  AOI22D1BWP U8411 ( .A1(vectorData2[137]), .A2(n5226), .B1(vectorData2[153]), 
        .B2(n5232), .ZN(n5178) );
  AO22D1BWP U8412 ( .A1(vectorData2[249]), .A2(n5229), .B1(vectorData2[41]), 
        .B2(n3601), .Z(n5180) );
  AOI22D1BWP U8413 ( .A1(vectorData2[73]), .A2(n5186), .B1(vectorData2[185]), 
        .B2(n5233), .ZN(n5182) );
  AOI22D1BWP U8414 ( .A1(n4681), .A2(vectorData2[9]), .B1(n4688), .B2(
        scalarData2[9]), .ZN(n3946) );
  ND4D1BWP U8415 ( .A1(n5246), .A2(n5245), .A3(n5244), .A4(n5243), .ZN(N4207)
         );
  AOI31D1BWP U8416 ( .A1(n5237), .A2(n5239), .A3(n5238), .B(n3661), .ZN(n5241)
         );
  AOI22D1BWP U8417 ( .A1(vectorData2[175]), .A2(n5230), .B1(vectorData2[255]), 
        .B2(n5229), .ZN(n5238) );
  AOI22D1BWP U8418 ( .A1(vectorData2[223]), .A2(n5228), .B1(vectorData2[207]), 
        .B2(n5227), .ZN(n5239) );
  OA211D1BWP U8419 ( .A1(n5236), .A2(n3673), .B(n5235), .C(n5234), .Z(n5237)
         );
  AOI22D1BWP U8420 ( .A1(vectorData2[191]), .A2(n5233), .B1(vectorData2[159]), 
        .B2(n5232), .ZN(n5234) );
  AOI22D1BWP U8421 ( .A1(vectorData2[127]), .A2(n5231), .B1(vectorData2[47]), 
        .B2(n3601), .ZN(n5235) );
  AOI22D1BWP U8422 ( .A1(vectorData2[15]), .A2(n4681), .B1(vectorData2[239]), 
        .B2(n4694), .ZN(n5242) );
  AOI22D1BWP U8423 ( .A1(scalarData2[15]), .A2(n4688), .B1(vectorData2[79]), 
        .B2(n4682), .ZN(n5244) );
  AOI22D1BWP U8424 ( .A1(vectorData2[95]), .A2(n4684), .B1(vectorData2[111]), 
        .B2(n4683), .ZN(n5245) );
  NR2XD0BWP U8425 ( .A1(n3672), .A2(n3661), .ZN(n4683) );
  AOI22D1BWP U8426 ( .A1(vectorData2[63]), .A2(n4686), .B1(vectorData2[31]), 
        .B2(n4685), .ZN(n5246) );
  OAI211D1BWP U8427 ( .A1(n128), .A2(n3670), .B(n4476), .C(n4475), .ZN(N4216)
         );
  ND3D1BWP U8428 ( .A1(n4478), .A2(n4474), .A3(result[0]), .ZN(n4475) );
  OAI222D1BWP U8429 ( .A1(n4699), .A2(n4539), .B1(n4538), .B2(n5277), .C1(
        n3670), .C2(n118), .ZN(N4226) );
  INVD1BWP U8430 ( .I(DataIn[10]), .ZN(n5277) );
  OAI222D1BWP U8431 ( .A1(\intadd_34/A[0] ), .A2(n4539), .B1(n4538), .B2(n5278), .C1(n3670), .C2(n117), .ZN(N4227) );
  OAI222D1BWP U8432 ( .A1(\intadd_34/A[1] ), .A2(n4539), .B1(n4538), .B2(n5279), .C1(n3670), .C2(n116), .ZN(N4228) );
  OAI222D1BWP U8433 ( .A1(\intadd_34/A[2] ), .A2(n4539), .B1(n4538), .B2(n5280), .C1(n3670), .C2(n115), .ZN(N4229) );
  OAI222D1BWP U8434 ( .A1(n3670), .A2(n114), .B1(n4538), .B2(n5281), .C1(n4539), .C2(\intadd_34/A[3] ), .ZN(N4230) );
  INVD1BWP U8435 ( .I(DataIn[14]), .ZN(n5281) );
  OAI222D1BWP U8436 ( .A1(n6037), .A2(n4539), .B1(n4538), .B2(n5283), .C1(
        n3670), .C2(n113), .ZN(N4231) );
  OAI222D1BWP U8437 ( .A1(n3670), .A2(n127), .B1(n4538), .B2(n5268), .C1(n4539), .C2(n4643), .ZN(N4217) );
  OAI222D1BWP U8438 ( .A1(n3670), .A2(n126), .B1(n4538), .B2(n5269), .C1(n4539), .C2(n4668), .ZN(N4218) );
  OAI222D1BWP U8439 ( .A1(n3670), .A2(n125), .B1(n4538), .B2(n5270), .C1(n4539), .C2(n6011), .ZN(N4219) );
  OAI222D1BWP U8440 ( .A1(n3670), .A2(n124), .B1(n4538), .B2(n5271), .C1(n4539), .C2(n4665), .ZN(N4220) );
  OAI222D1BWP U8441 ( .A1(n3670), .A2(n123), .B1(n4539), .B2(n4664), .C1(n4538), .C2(n5272), .ZN(N4221) );
  OAI222D1BWP U8442 ( .A1(n3670), .A2(n122), .B1(n4539), .B2(n4661), .C1(n4538), .C2(n5273), .ZN(N4222) );
  OAI222D1BWP U8443 ( .A1(n3670), .A2(n121), .B1(n4539), .B2(n4655), .C1(n4538), .C2(n5274), .ZN(N4223) );
  OAI222D1BWP U8444 ( .A1(n3670), .A2(n120), .B1(n4539), .B2(n4652), .C1(n4538), .C2(n5275), .ZN(N4224) );
  OAI222D1BWP U8445 ( .A1(n3670), .A2(n119), .B1(n4539), .B2(n4651), .C1(n4538), .C2(n5276), .ZN(N4225) );
  OAI31D1BWP U8446 ( .A1(cycles[4]), .A2(n5298), .A3(n5302), .B(n5249), .ZN(
        n5250) );
  OAI22D1BWP U8447 ( .A1(n4967), .A2(n4918), .B1(n4917), .B2(n4962), .ZN(N1820) );
  OAI32D1BWP U8448 ( .A1(n4700), .A2(n4956), .A3(n4916), .B1(n4915), .B2(n4955), .ZN(n4917) );
  NR2XD0BWP U8449 ( .A1(n4963), .A2(n4942), .ZN(n4916) );
  NR2XD0BWP U8450 ( .A1(n5249), .A2(result[10]), .ZN(n4918) );
  OAI21D1BWP U8451 ( .A1(n4467), .A2(n4557), .B(n4466), .ZN(N4212) );
  OAI21D1BWP U8452 ( .A1(n4467), .A2(n4560), .B(n4466), .ZN(N4213) );
  NR2XD0BWP U8453 ( .A1(n6040), .A2(n5248), .ZN(n4467) );
  AO211D1BWP U8454 ( .A1(n4073), .A2(scalarData1[13]), .B(n3938), .C(n3937), 
        .Z(N4189) );
  AO22D1BWP U8455 ( .A1(n4072), .A2(vectorData1[13]), .B1(n4071), .B2(Addr[13]), .Z(n3937) );
  ND4D1BWP U8456 ( .A1(n7159), .A2(n7160), .A3(n7161), .A4(n7162), .ZN(
        vectorData1[13]) );
  AOI22D1BWP U8457 ( .A1(n3576), .A2(\vrf/regTable[5][13] ), .B1(n3567), .B2(
        \vrf/regTable[7][13] ), .ZN(n7162) );
  AOI22D1BWP U8458 ( .A1(n3574), .A2(\vrf/regTable[4][13] ), .B1(n3570), .B2(
        \vrf/regTable[6][13] ), .ZN(n7161) );
  AOI22D1BWP U8459 ( .A1(n3579), .A2(\vrf/regTable[1][13] ), .B1(n3575), .B2(
        \vrf/regTable[3][13] ), .ZN(n7160) );
  AOI22D1BWP U8460 ( .A1(n3581), .A2(\vrf/regTable[0][13] ), .B1(n3572), .B2(
        \vrf/regTable[2][13] ), .ZN(n7159) );
  AOI31D1BWP U8461 ( .A1(n5110), .A2(n5109), .A3(n5111), .B(n4070), .ZN(n3938)
         );
  NR2XD0BWP U8462 ( .A1(n3732), .A2(n4394), .ZN(n4695) );
  AOI22D1BWP U8463 ( .A1(n5185), .A2(vectorData1[93]), .B1(n5186), .B2(
        vectorData1[77]), .ZN(n5111) );
  ND4D1BWP U8464 ( .A1(n7411), .A2(n7412), .A3(n7413), .A4(n7414), .ZN(
        vectorData1[77]) );
  AOI22D1BWP U8465 ( .A1(n3576), .A2(\vrf/regTable[5][77] ), .B1(n3595), .B2(
        \vrf/regTable[7][77] ), .ZN(n7414) );
  AOI22D1BWP U8466 ( .A1(n3574), .A2(\vrf/regTable[4][77] ), .B1(n3596), .B2(
        \vrf/regTable[6][77] ), .ZN(n7413) );
  AOI22D1BWP U8467 ( .A1(n3579), .A2(\vrf/regTable[1][77] ), .B1(n3599), .B2(
        \vrf/regTable[3][77] ), .ZN(n7412) );
  AOI22D1BWP U8468 ( .A1(n3581), .A2(\vrf/regTable[0][77] ), .B1(n3594), .B2(
        \vrf/regTable[2][77] ), .ZN(n7411) );
  ND4D1BWP U8469 ( .A1(n7475), .A2(n7476), .A3(n7477), .A4(n7478), .ZN(
        vectorData1[93]) );
  AOI22D1BWP U8470 ( .A1(n3576), .A2(\vrf/regTable[5][93] ), .B1(n3567), .B2(
        \vrf/regTable[7][93] ), .ZN(n7478) );
  AOI22D1BWP U8471 ( .A1(n3574), .A2(\vrf/regTable[4][93] ), .B1(n3570), .B2(
        \vrf/regTable[6][93] ), .ZN(n7477) );
  AOI22D1BWP U8472 ( .A1(n3579), .A2(\vrf/regTable[1][93] ), .B1(n3575), .B2(
        \vrf/regTable[3][93] ), .ZN(n7476) );
  AOI22D1BWP U8473 ( .A1(n3581), .A2(\vrf/regTable[0][93] ), .B1(n3572), .B2(
        \vrf/regTable[2][93] ), .ZN(n7475) );
  AOI211XD0BWP U8474 ( .A1(n5187), .A2(vectorData1[237]), .B(n5108), .C(n5107), 
        .ZN(n5109) );
  ND4D1BWP U8475 ( .A1(n5106), .A2(n5105), .A3(n5104), .A4(n5103), .ZN(n5107)
         );
  AOI22D1BWP U8476 ( .A1(n5229), .A2(vectorData1[253]), .B1(n5227), .B2(
        vectorData1[205]), .ZN(n5103) );
  ND4D1BWP U8477 ( .A1(n7923), .A2(n7924), .A3(n7925), .A4(n7926), .ZN(
        vectorData1[205]) );
  AOI22D1BWP U8478 ( .A1(n3576), .A2(\vrf/regTable[5][205] ), .B1(n7118), .B2(
        \vrf/regTable[7][205] ), .ZN(n7926) );
  AOI22D1BWP U8479 ( .A1(n3574), .A2(\vrf/regTable[4][205] ), .B1(n7116), .B2(
        \vrf/regTable[6][205] ), .ZN(n7925) );
  AOI22D1BWP U8480 ( .A1(n3579), .A2(\vrf/regTable[1][205] ), .B1(n7114), .B2(
        \vrf/regTable[3][205] ), .ZN(n7924) );
  AOI22D1BWP U8481 ( .A1(n3581), .A2(\vrf/regTable[0][205] ), .B1(n7110), .B2(
        \vrf/regTable[2][205] ), .ZN(n7923) );
  ND4D1BWP U8482 ( .A1(n8115), .A2(n8116), .A3(n8117), .A4(n8118), .ZN(
        vectorData1[253]) );
  AOI22D1BWP U8483 ( .A1(n3576), .A2(\vrf/regTable[5][253] ), .B1(n3595), .B2(
        \vrf/regTable[7][253] ), .ZN(n8118) );
  AOI22D1BWP U8484 ( .A1(n3574), .A2(\vrf/regTable[4][253] ), .B1(n3596), .B2(
        \vrf/regTable[6][253] ), .ZN(n8117) );
  AOI22D1BWP U8485 ( .A1(n3579), .A2(\vrf/regTable[1][253] ), .B1(n3599), .B2(
        \vrf/regTable[3][253] ), .ZN(n8116) );
  AOI22D1BWP U8486 ( .A1(n3581), .A2(\vrf/regTable[0][253] ), .B1(n3594), .B2(
        \vrf/regTable[2][253] ), .ZN(n8115) );
  AOI22D1BWP U8487 ( .A1(n5226), .A2(vectorData1[141]), .B1(n5231), .B2(
        vectorData1[125]), .ZN(n5104) );
  ND4D1BWP U8488 ( .A1(n7603), .A2(n7604), .A3(n7605), .A4(n7606), .ZN(
        vectorData1[125]) );
  AOI22D1BWP U8489 ( .A1(n3576), .A2(\vrf/regTable[5][125] ), .B1(n3567), .B2(
        \vrf/regTable[7][125] ), .ZN(n7606) );
  AOI22D1BWP U8490 ( .A1(n3574), .A2(\vrf/regTable[4][125] ), .B1(n3570), .B2(
        \vrf/regTable[6][125] ), .ZN(n7605) );
  AOI22D1BWP U8491 ( .A1(n3579), .A2(\vrf/regTable[1][125] ), .B1(n3575), .B2(
        \vrf/regTable[3][125] ), .ZN(n7604) );
  AOI22D1BWP U8492 ( .A1(n3581), .A2(\vrf/regTable[0][125] ), .B1(n3572), .B2(
        \vrf/regTable[2][125] ), .ZN(n7603) );
  ND4D1BWP U8493 ( .A1(n7667), .A2(n7668), .A3(n7669), .A4(n7670), .ZN(
        vectorData1[141]) );
  AOI22D1BWP U8494 ( .A1(n3576), .A2(\vrf/regTable[5][141] ), .B1(n3567), .B2(
        \vrf/regTable[7][141] ), .ZN(n7670) );
  AOI22D1BWP U8495 ( .A1(n3574), .A2(\vrf/regTable[4][141] ), .B1(n3570), .B2(
        \vrf/regTable[6][141] ), .ZN(n7669) );
  AOI22D1BWP U8496 ( .A1(n3579), .A2(\vrf/regTable[1][141] ), .B1(n3599), .B2(
        \vrf/regTable[3][141] ), .ZN(n7668) );
  AOI22D1BWP U8497 ( .A1(n3581), .A2(\vrf/regTable[0][141] ), .B1(n3572), .B2(
        \vrf/regTable[2][141] ), .ZN(n7667) );
  AOI22D1BWP U8498 ( .A1(n5213), .A2(vectorData1[109]), .B1(n5232), .B2(
        vectorData1[157]), .ZN(n5105) );
  ND4D1BWP U8499 ( .A1(n7731), .A2(n7732), .A3(n7733), .A4(n7734), .ZN(
        vectorData1[157]) );
  AOI22D1BWP U8500 ( .A1(n3576), .A2(\vrf/regTable[5][157] ), .B1(n3595), .B2(
        \vrf/regTable[7][157] ), .ZN(n7734) );
  AOI22D1BWP U8501 ( .A1(n3574), .A2(\vrf/regTable[4][157] ), .B1(n3596), .B2(
        \vrf/regTable[6][157] ), .ZN(n7733) );
  AOI22D1BWP U8502 ( .A1(n3579), .A2(\vrf/regTable[1][157] ), .B1(n3575), .B2(
        \vrf/regTable[3][157] ), .ZN(n7732) );
  AOI22D1BWP U8503 ( .A1(n3581), .A2(\vrf/regTable[0][157] ), .B1(n3594), .B2(
        \vrf/regTable[2][157] ), .ZN(n7731) );
  ND4D1BWP U8504 ( .A1(n7539), .A2(n7540), .A3(n7541), .A4(n7542), .ZN(
        vectorData1[109]) );
  AOI22D1BWP U8505 ( .A1(n3576), .A2(\vrf/regTable[5][109] ), .B1(n3595), .B2(
        \vrf/regTable[7][109] ), .ZN(n7542) );
  AOI22D1BWP U8506 ( .A1(n3574), .A2(\vrf/regTable[4][109] ), .B1(n3596), .B2(
        \vrf/regTable[6][109] ), .ZN(n7541) );
  AOI22D1BWP U8507 ( .A1(n3579), .A2(\vrf/regTable[1][109] ), .B1(n3599), .B2(
        \vrf/regTable[3][109] ), .ZN(n7540) );
  AOI22D1BWP U8508 ( .A1(n3581), .A2(\vrf/regTable[0][109] ), .B1(n3594), .B2(
        \vrf/regTable[2][109] ), .ZN(n7539) );
  AOI22D1BWP U8509 ( .A1(n5233), .A2(vectorData1[189]), .B1(n5184), .B2(
        vectorData1[29]), .ZN(n5106) );
  ND4D1BWP U8510 ( .A1(n7219), .A2(n7220), .A3(n7221), .A4(n7222), .ZN(
        vectorData1[29]) );
  AOI22D1BWP U8511 ( .A1(n3576), .A2(\vrf/regTable[5][29] ), .B1(n3595), .B2(
        \vrf/regTable[7][29] ), .ZN(n7222) );
  AOI22D1BWP U8512 ( .A1(n3574), .A2(\vrf/regTable[4][29] ), .B1(n3596), .B2(
        \vrf/regTable[6][29] ), .ZN(n7221) );
  AOI22D1BWP U8513 ( .A1(n3579), .A2(\vrf/regTable[1][29] ), .B1(n3599), .B2(
        \vrf/regTable[3][29] ), .ZN(n7220) );
  AOI22D1BWP U8514 ( .A1(n3581), .A2(\vrf/regTable[0][29] ), .B1(n3594), .B2(
        \vrf/regTable[2][29] ), .ZN(n7219) );
  ND4D1BWP U8515 ( .A1(n7859), .A2(n7860), .A3(n7861), .A4(n7862), .ZN(
        vectorData1[189]) );
  AOI22D1BWP U8516 ( .A1(n3576), .A2(\vrf/regTable[5][189] ), .B1(n3567), .B2(
        \vrf/regTable[7][189] ), .ZN(n7862) );
  AOI22D1BWP U8517 ( .A1(n3574), .A2(\vrf/regTable[4][189] ), .B1(n3570), .B2(
        \vrf/regTable[6][189] ), .ZN(n7861) );
  AOI22D1BWP U8518 ( .A1(n3579), .A2(\vrf/regTable[1][189] ), .B1(n3575), .B2(
        \vrf/regTable[3][189] ), .ZN(n7860) );
  AOI22D1BWP U8519 ( .A1(n3581), .A2(\vrf/regTable[0][189] ), .B1(n3572), .B2(
        \vrf/regTable[2][189] ), .ZN(n7859) );
  AO22D1BWP U8520 ( .A1(n5188), .A2(vectorData1[61]), .B1(n5230), .B2(
        vectorData1[173]), .Z(n5108) );
  ND4D1BWP U8521 ( .A1(n7795), .A2(n7796), .A3(n7797), .A4(n7798), .ZN(
        vectorData1[173]) );
  AOI22D1BWP U8522 ( .A1(n3576), .A2(\vrf/regTable[5][173] ), .B1(n7118), .B2(
        \vrf/regTable[7][173] ), .ZN(n7798) );
  AOI22D1BWP U8523 ( .A1(n3574), .A2(\vrf/regTable[4][173] ), .B1(n7116), .B2(
        \vrf/regTable[6][173] ), .ZN(n7797) );
  AOI22D1BWP U8524 ( .A1(n3579), .A2(\vrf/regTable[1][173] ), .B1(n7114), .B2(
        \vrf/regTable[3][173] ), .ZN(n7796) );
  AOI22D1BWP U8525 ( .A1(n3581), .A2(\vrf/regTable[0][173] ), .B1(n7110), .B2(
        \vrf/regTable[2][173] ), .ZN(n7795) );
  ND4D1BWP U8526 ( .A1(n7347), .A2(n7348), .A3(n7349), .A4(n7350), .ZN(
        vectorData1[61]) );
  AOI22D1BWP U8527 ( .A1(n3576), .A2(\vrf/regTable[5][61] ), .B1(n3567), .B2(
        \vrf/regTable[7][61] ), .ZN(n7350) );
  AOI22D1BWP U8528 ( .A1(n3574), .A2(\vrf/regTable[4][61] ), .B1(n3570), .B2(
        \vrf/regTable[6][61] ), .ZN(n7349) );
  AOI22D1BWP U8529 ( .A1(n3579), .A2(\vrf/regTable[1][61] ), .B1(n3575), .B2(
        \vrf/regTable[3][61] ), .ZN(n7348) );
  AOI22D1BWP U8530 ( .A1(n3581), .A2(\vrf/regTable[0][61] ), .B1(n3572), .B2(
        \vrf/regTable[2][61] ), .ZN(n7347) );
  ND4D1BWP U8531 ( .A1(n8051), .A2(n8052), .A3(n8053), .A4(n8054), .ZN(
        vectorData1[237]) );
  AOI22D1BWP U8532 ( .A1(n3576), .A2(\vrf/regTable[5][237] ), .B1(n3595), .B2(
        \vrf/regTable[7][237] ), .ZN(n8054) );
  AOI22D1BWP U8533 ( .A1(n3574), .A2(\vrf/regTable[4][237] ), .B1(n3596), .B2(
        \vrf/regTable[6][237] ), .ZN(n8053) );
  AOI22D1BWP U8534 ( .A1(n3579), .A2(\vrf/regTable[1][237] ), .B1(n3599), .B2(
        \vrf/regTable[3][237] ), .ZN(n8052) );
  AOI22D1BWP U8535 ( .A1(n3581), .A2(\vrf/regTable[0][237] ), .B1(n3594), .B2(
        \vrf/regTable[2][237] ), .ZN(n8051) );
  AOI22D1BWP U8536 ( .A1(n5228), .A2(vectorData1[221]), .B1(n3601), .B2(
        vectorData1[45]), .ZN(n5110) );
  ND4D1BWP U8537 ( .A1(n7283), .A2(n7284), .A3(n7285), .A4(n7286), .ZN(
        vectorData1[45]) );
  AOI22D1BWP U8538 ( .A1(n3576), .A2(\vrf/regTable[5][45] ), .B1(n3595), .B2(
        \vrf/regTable[7][45] ), .ZN(n7286) );
  AOI22D1BWP U8539 ( .A1(n3574), .A2(\vrf/regTable[4][45] ), .B1(n3596), .B2(
        \vrf/regTable[6][45] ), .ZN(n7285) );
  AOI22D1BWP U8540 ( .A1(n3579), .A2(\vrf/regTable[1][45] ), .B1(n3599), .B2(
        \vrf/regTable[3][45] ), .ZN(n7284) );
  AOI22D1BWP U8541 ( .A1(n3581), .A2(\vrf/regTable[0][45] ), .B1(n3594), .B2(
        \vrf/regTable[2][45] ), .ZN(n7283) );
  ND4D1BWP U8542 ( .A1(n7987), .A2(n7988), .A3(n7989), .A4(n7990), .ZN(
        vectorData1[221]) );
  AOI22D1BWP U8543 ( .A1(n3576), .A2(\vrf/regTable[5][221] ), .B1(n3595), .B2(
        \vrf/regTable[7][221] ), .ZN(n7990) );
  NR2XD0BWP U8544 ( .A1(n7113), .A2(n4619), .ZN(n7118) );
  NR2XD0BWP U8545 ( .A1(n7111), .A2(n4619), .ZN(n7117) );
  AOI22D1BWP U8546 ( .A1(n3574), .A2(\vrf/regTable[4][221] ), .B1(n3596), .B2(
        \vrf/regTable[6][221] ), .ZN(n7989) );
  NR2XD0BWP U8547 ( .A1(n7109), .A2(n4619), .ZN(n7116) );
  AOI22D1BWP U8548 ( .A1(n3579), .A2(\vrf/regTable[1][221] ), .B1(n3599), .B2(
        \vrf/regTable[3][221] ), .ZN(n7988) );
  NR2XD0BWP U8549 ( .A1(n7113), .A2(\vrf/N11 ), .ZN(n7114) );
  NR2XD0BWP U8550 ( .A1(n7111), .A2(\vrf/N11 ), .ZN(n7112) );
  AOI22D1BWP U8551 ( .A1(n3581), .A2(\vrf/regTable[0][221] ), .B1(n3594), .B2(
        \vrf/regTable[2][221] ), .ZN(n7987) );
  NR2XD0BWP U8552 ( .A1(n7109), .A2(\vrf/N11 ), .ZN(n7110) );
  ND4D1BWP U8553 ( .A1(n8329), .A2(n8330), .A3(n8331), .A4(n8332), .ZN(
        scalarData1[13]) );
  AOI22D1BWP U8554 ( .A1(n8287), .A2(\srf/regTable[5][13] ), .B1(n8288), .B2(
        \srf/regTable[7][13] ), .ZN(n8332) );
  NR2XD0BWP U8555 ( .A1(n8283), .A2(n4619), .ZN(n8288) );
  NR2XD0BWP U8556 ( .A1(n8281), .A2(n4619), .ZN(n8287) );
  AOI22D1BWP U8557 ( .A1(n8285), .A2(\srf/regTable[4][13] ), .B1(n8286), .B2(
        \srf/regTable[6][13] ), .ZN(n8331) );
  NR2XD0BWP U8558 ( .A1(n8279), .A2(n4619), .ZN(n8286) );
  AOI22D1BWP U8559 ( .A1(n8282), .A2(\srf/regTable[1][13] ), .B1(n8284), .B2(
        \srf/regTable[3][13] ), .ZN(n8330) );
  NR2XD0BWP U8560 ( .A1(n8283), .A2(\vrf/N11 ), .ZN(n8284) );
  NR2XD0BWP U8561 ( .A1(n8281), .A2(\vrf/N11 ), .ZN(n8282) );
  AOI22D1BWP U8562 ( .A1(n8278), .A2(\srf/regTable[0][13] ), .B1(n8280), .B2(
        \srf/regTable[2][13] ), .ZN(n8329) );
  NR2XD0BWP U8563 ( .A1(n8279), .A2(\vrf/N11 ), .ZN(n8280) );
  OAI22D1BWP U8564 ( .A1(n4561), .A2(n4560), .B1(n4559), .B2(n4558), .ZN(
        \vrf/N10 ) );
  OAI22D1BWP U8565 ( .A1(n4561), .A2(n4557), .B1(n4556), .B2(n4558), .ZN(
        \vrf/N9 ) );
  OAI22D1BWP U8566 ( .A1(n4967), .A2(n4959), .B1(n4960), .B2(n4962), .ZN(N1823) );
  AOI222D1BWP U8567 ( .A1(n4958), .A2(n4961), .B1(n4957), .B2(n4956), .C1(
        n4955), .C2(n4954), .ZN(n4960) );
  IND3D1BWP U8568 ( .A1(n4952), .B1(n4951), .B2(n4950), .ZN(n4958) );
  OAI211D1BWP U8569 ( .A1(n4957), .A2(n4949), .B(n4948), .C(n4947), .ZN(n4950)
         );
  AOI22D1BWP U8570 ( .A1(n4951), .A2(n4952), .B1(n4387), .B2(n4946), .ZN(n4949) );
  MAOI222D1BWP U8571 ( .A(n4945), .B(n4944), .C(n4943), .ZN(n4946) );
  AOI32D1BWP U8572 ( .A1(n4941), .A2(n4940), .A3(n4939), .B1(n4938), .B2(n4940), .ZN(n4944) );
  OAI21D1BWP U8573 ( .A1(n4937), .A2(n4936), .B(n4935), .ZN(n4939) );
  NR2XD0BWP U8574 ( .A1(n4938), .A2(n4933), .ZN(n4951) );
  XNR2D1BWP U8575 ( .A1(n4905), .A2(n4869), .ZN(n4931) );
  XNR2D1BWP U8576 ( .A1(n4908), .A2(n4907), .ZN(n4932) );
  INR2D1BWP U8577 ( .A1(n4905), .B1(n4904), .ZN(n4908) );
  INR2D1BWP U8578 ( .A1(n4930), .B1(n4929), .ZN(n4935) );
  OAI21D1BWP U8579 ( .A1(n4903), .A2(n4353), .B(n4354), .ZN(n4155) );
  INR2D1BWP U8580 ( .A1(n4928), .B1(n4927), .ZN(n4941) );
  OAI31D1BWP U8581 ( .A1(n4899), .A2(n4898), .A3(n4903), .B(n4897), .ZN(n4914)
         );
  OAI21D1BWP U8582 ( .A1(n4903), .A2(n4898), .B(n4899), .ZN(n4897) );
  OAI31D1BWP U8583 ( .A1(n4902), .A2(n4901), .A3(n4903), .B(n4900), .ZN(n4928)
         );
  OAI21D1BWP U8584 ( .A1(n4903), .A2(n4901), .B(n4902), .ZN(n4900) );
  NR2XD0BWP U8585 ( .A1(n5249), .A2(result[13]), .ZN(n4959) );
  OAI22D1BWP U8586 ( .A1(n4820), .A2(n4810), .B1(n4816), .B2(n4811), .ZN(
        \mult_x_153/n152 ) );
  OAI22D1BWP U8587 ( .A1(n5554), .A2(n4794), .B1(n4793), .B2(n4797), .ZN(
        \mult_x_153/n132 ) );
  AOI22D1BWP U8588 ( .A1(op1[9]), .A2(n4670), .B1(op2[2]), .B2(n3680), .ZN(
        n4797) );
  OAI32D1BWP U8589 ( .A1(\mult_x_153/n98 ), .A2(\mult_x_153/n148 ), .A3(
        \mult_x_153/n136 ), .B1(n4786), .B2(\mult_x_153/n98 ), .ZN(
        \mult_x_153/n99 ) );
  OAI22D1BWP U8590 ( .A1(n5576), .A2(n4826), .B1(n4856), .B2(n5562), .ZN(
        \mult_x_153/n170 ) );
  OAI22D1BWP U8591 ( .A1(n4967), .A2(n4921), .B1(n4920), .B2(n4962), .ZN(N1821) );
  AOI211XD0BWP U8592 ( .A1(n4956), .A2(n4945), .B(n4919), .C(n4924), .ZN(n4920) );
  IND2D1BWP U8593 ( .A1(n4936), .B1(n4937), .ZN(n4948) );
  MUX2ND0BWP U8594 ( .I0(n4868), .I1(n4165), .S(n4903), .ZN(n4937) );
  MUX2ND0BWP U8595 ( .I0(n4161), .I1(n4160), .S(n4903), .ZN(n4913) );
  OAI31D1BWP U8596 ( .A1(n4903), .A2(n4894), .A3(n4895), .B(n4893), .ZN(n4912)
         );
  OAI21D1BWP U8597 ( .A1(n4903), .A2(n4894), .B(n4895), .ZN(n4893) );
  NR2XD0BWP U8598 ( .A1(n4961), .A2(n4955), .ZN(n4956) );
  ND3D1BWP U8599 ( .A1(n4146), .A2(n4338), .A3(n4100), .ZN(n4966) );
  NR2XD0BWP U8600 ( .A1(n5249), .A2(result[11]), .ZN(n4921) );
  OA211D1BWP U8601 ( .A1(n4076), .A2(n4075), .B(n5249), .C(n4074), .Z(n4639)
         );
  ND3D1BWP U8602 ( .A1(scalarToLoad[10]), .A2(scalarToLoad[14]), .A3(
        scalarToLoad[13]), .ZN(n4075) );
  XNR2D1BWP U8603 ( .A1(n4389), .A2(n4388), .ZN(n4632) );
  NR2XD0BWP U8604 ( .A1(n4882), .A2(n4633), .ZN(n4388) );
  XOR2D1BWP U8605 ( .A1(n4889), .A2(n4879), .Z(n4934) );
  NR2XD0BWP U8606 ( .A1(n4870), .A2(n4903), .ZN(n4905) );
  NR2XD0BWP U8607 ( .A1(n4915), .A2(n4945), .ZN(n4881) );
  XOR2D1BWP U8608 ( .A1(n4891), .A2(n4880), .Z(n4945) );
  MUX2ND0BWP U8609 ( .I0(n4633), .I1(n4957), .S(n4964), .ZN(n4953) );
  NR2XD0BWP U8610 ( .A1(n4700), .A2(n4891), .ZN(n4922) );
  XOR2D1BWP U8611 ( .A1(n4878), .A2(n4890), .Z(n4915) );
  XOR2D1BWP U8612 ( .A1(n4633), .A2(n4882), .Z(n4957) );
  NR2XD0BWP U8613 ( .A1(n4880), .A2(n4891), .ZN(n4879) );
  NR2XD0BWP U8614 ( .A1(n4888), .A2(n4903), .ZN(n4878) );
  ND3D1BWP U8615 ( .A1(n4386), .A2(n4385), .A3(n4390), .ZN(n4903) );
  ND4D1BWP U8616 ( .A1(n4360), .A2(n4382), .A3(n4121), .A4(n4362), .ZN(n4390)
         );
  NR2XD0BWP U8617 ( .A1(n4635), .A2(n4884), .ZN(n4121) );
  AOI21D1BWP U8618 ( .A1(n4884), .A2(n4379), .B(n4378), .ZN(n4633) );
  OAI22D1BWP U8619 ( .A1(n4379), .A2(n4377), .B1(n4867), .B2(n4887), .ZN(n4378) );
  NR2XD0BWP U8620 ( .A1(n4877), .A2(n4374), .ZN(n4379) );
  ND3D1BWP U8621 ( .A1(n4164), .A2(n4139), .A3(n4116), .ZN(n4386) );
  NR4D0BWP U8622 ( .A1(N1463), .A2(N1462), .A3(N1460), .A4(N1458), .ZN(n4112)
         );
  NR4D0BWP U8623 ( .A1(N1467), .A2(N1466), .A3(N1465), .A4(N1464), .ZN(n4113)
         );
  AOI211XD0BWP U8624 ( .A1(N1457), .A2(n4374), .B(N1468), .C(N1469), .ZN(n4114) );
  AOI211XD0BWP U8625 ( .A1(N1470), .A2(N1483), .B(N1461), .C(N1459), .ZN(n4115) );
  AO211D1BWP U8626 ( .A1(n4373), .A2(n4876), .B(n4372), .C(n4371), .Z(n4889)
         );
  OAI22D1BWP U8627 ( .A1(n4635), .A2(n4370), .B1(n4876), .B2(n4369), .ZN(n4371) );
  OA211D1BWP U8628 ( .A1(n4368), .A2(n4367), .B(N1483), .C(n4877), .Z(n4372)
         );
  AOI21D1BWP U8629 ( .A1(n4875), .A2(n4635), .B(n4874), .ZN(n4876) );
  AOI211XD0BWP U8630 ( .A1(n4384), .A2(n4383), .B(n4382), .C(n4381), .ZN(n4389) );
  NR2XD0BWP U8631 ( .A1(n4887), .A2(n4380), .ZN(n4381) );
  XNR2D1BWP U8632 ( .A1(n4885), .A2(n4383), .ZN(n4380) );
  NR2XD0BWP U8633 ( .A1(n4635), .A2(n4875), .ZN(n4874) );
  AOI31D1BWP U8634 ( .A1(n4119), .A2(n4383), .A3(n4375), .B(n4118), .ZN(n4382)
         );
  OAI21D1BWP U8635 ( .A1(n4884), .A2(n4877), .B(n4886), .ZN(n4863) );
  MUX2ND0BWP U8636 ( .I0(result[13]), .I1(scalarToLoad[13]), .S(\intadd_34/CO ), .ZN(n4884) );
  MUX2ND0BWP U8637 ( .I0(result[12]), .I1(scalarToLoad[12]), .S(\intadd_34/n1 ), .ZN(n4635) );
  NR2XD0BWP U8638 ( .A1(n4120), .A2(n4360), .ZN(n4368) );
  NR2XD0BWP U8639 ( .A1(result[14]), .A2(scalarToLoad[14]), .ZN(n4886) );
  OAI21D1BWP U8640 ( .A1(n4360), .A2(n4357), .B(n4356), .ZN(n4890) );
  AOI21D1BWP U8641 ( .A1(n4355), .A2(n4366), .B(n4384), .ZN(n4357) );
  OAI211D1BWP U8642 ( .A1(n4153), .A2(n4148), .B(n4105), .C(n4104), .ZN(n4907)
         );
  OA211D1BWP U8643 ( .A1(n4123), .A2(n4345), .B(n4099), .C(n4098), .Z(n4105)
         );
  AOI22D1BWP U8644 ( .A1(N1480), .A2(n4341), .B1(N1483), .B2(N1481), .ZN(n4099) );
  ND4D1BWP U8645 ( .A1(n4132), .A2(n4131), .A3(n4130), .A4(n4129), .ZN(n4872)
         );
  ND3D1BWP U8646 ( .A1(n4143), .A2(n4349), .A3(n4142), .ZN(n4129) );
  MUX2ND0BWP U8647 ( .I0(N1477), .I1(N1478), .S(n4355), .ZN(n4123) );
  AOI22D1BWP U8648 ( .A1(N1479), .A2(N1483), .B1(N1478), .B2(n4341), .ZN(n4132) );
  NR2XD0BWP U8649 ( .A1(n4898), .A2(n4899), .ZN(n4873) );
  AOI211XD0BWP U8650 ( .A1(n4151), .A2(n4373), .B(n4111), .C(n4110), .ZN(n4904) );
  OAI22D1BWP U8651 ( .A1(n4340), .A2(n4345), .B1(n4149), .B2(n4109), .ZN(n4110) );
  OAI21D1BWP U8652 ( .A1(n4346), .A2(n4122), .B(n4108), .ZN(n4111) );
  AOI22D1BWP U8653 ( .A1(N1480), .A2(N1483), .B1(N1479), .B2(n4341), .ZN(n4108) );
  IOA21D1BWP U8654 ( .A1(n4373), .A2(n4865), .B(n4350), .ZN(n4871) );
  AOI21D1BWP U8655 ( .A1(n4349), .A2(n4348), .B(n4347), .ZN(n4350) );
  OAI211D1BWP U8656 ( .A1(n4346), .A2(n4345), .B(n4344), .C(n4343), .ZN(n4347)
         );
  AOI22D1BWP U8657 ( .A1(N1483), .A2(N1482), .B1(N1481), .B2(n4341), .ZN(n4344) );
  NR2XD0BWP U8658 ( .A1(n4100), .A2(n4376), .ZN(n4349) );
  OAI21D1BWP U8659 ( .A1(n4159), .A2(n4160), .B(n4894), .ZN(n4892) );
  AOI21D1BWP U8660 ( .A1(n4636), .A2(n4865), .B(n4864), .ZN(n4899) );
  AO222D1BWP U8661 ( .A1(n4341), .A2(N1477), .B1(N1478), .B2(N1483), .C1(n4373), .C2(n4348), .Z(n4864) );
  MUX2ND0BWP U8662 ( .I0(n4340), .I1(n4339), .S(n4359), .ZN(n4865) );
  MUX2ND0BWP U8663 ( .I0(N1476), .I1(N1477), .S(n4355), .ZN(n4340) );
  XOR2D1BWP U8664 ( .A1(n4164), .A2(n4163), .Z(n4868) );
  MUX2ND0BWP U8665 ( .I0(n4124), .I1(n4126), .S(n4359), .ZN(n4153) );
  NR2XD0BWP U8666 ( .A1(n4353), .A2(n4354), .ZN(n4634) );
  OAI31D1BWP U8667 ( .A1(n4146), .A2(n4145), .A3(n4376), .B(n4144), .ZN(n4895)
         );
  AOI22D1BWP U8668 ( .A1(N1483), .A2(N1475), .B1(N1474), .B2(n4341), .ZN(n4144) );
  AOI22D1BWP U8669 ( .A1(n4143), .A2(n4142), .B1(n4141), .B2(n4866), .ZN(n4145) );
  MUX2ND0BWP U8670 ( .I0(n4128), .I1(n4127), .S(n4359), .ZN(n4141) );
  MUX2ND0BWP U8671 ( .I0(n4092), .I1(n4091), .S(n4355), .ZN(n4126) );
  AO222D1BWP U8672 ( .A1(n4341), .A2(N1473), .B1(N1483), .B2(N1474), .C1(n4636), .C2(n4348), .Z(n4160) );
  MUX2ND0BWP U8673 ( .I0(n4140), .I1(n4149), .S(n4359), .ZN(n4348) );
  NR2XD0BWP U8674 ( .A1(n4163), .A2(n4164), .ZN(n4159) );
  AOI222D1BWP U8675 ( .A1(N1473), .A2(N1483), .B1(N1472), .B2(n4384), .C1(
        n4636), .C2(n4152), .ZN(n4164) );
  MUX2ND0BWP U8676 ( .I0(n4127), .I1(n4103), .S(n4359), .ZN(n4152) );
  MUX2ND0BWP U8677 ( .I0(N1471), .I1(N1472), .S(n4355), .ZN(n4127) );
  IND3D1BWP U8678 ( .A1(n4139), .B1(n4138), .B2(n4385), .ZN(n4163) );
  OAI21D1BWP U8679 ( .A1(n4149), .A2(n4122), .B(n4117), .ZN(n4385) );
  AOI22D1BWP U8680 ( .A1(N1472), .A2(N1483), .B1(N1471), .B2(n4341), .ZN(n4117) );
  NR4D0BWP U8681 ( .A1(n4137), .A2(n4136), .A3(n4135), .A4(n4134), .ZN(n4138)
         );
  ND4D1BWP U8682 ( .A1(N1463), .A2(N1462), .A3(N1460), .A4(N1458), .ZN(n4134)
         );
  XOR2D1BWP U8683 ( .A1(\DP_OP_487J11_125_9213/n26 ), .A2(
        \DP_OP_487J11_125_9213/n55 ), .Z(N1458) );
  XOR2D1BWP U8684 ( .A1(\DP_OP_487J11_125_9213/n24 ), .A2(
        \DP_OP_487J11_125_9213/n53 ), .Z(N1460) );
  XOR2D1BWP U8685 ( .A1(\DP_OP_487J11_125_9213/n22 ), .A2(
        \DP_OP_487J11_125_9213/n51 ), .Z(N1462) );
  XOR2D1BWP U8686 ( .A1(\DP_OP_487J11_125_9213/n21 ), .A2(
        \DP_OP_487J11_125_9213/n50 ), .Z(N1463) );
  ND4D1BWP U8687 ( .A1(N1467), .A2(N1466), .A3(N1465), .A4(N1464), .ZN(n4135)
         );
  XOR2D1BWP U8688 ( .A1(\DP_OP_487J11_125_9213/n20 ), .A2(
        \DP_OP_487J11_125_9213/n49 ), .Z(N1464) );
  XOR2D1BWP U8689 ( .A1(\DP_OP_487J11_125_9213/n19 ), .A2(
        \DP_OP_487J11_125_9213/n48 ), .Z(N1465) );
  XOR2D1BWP U8690 ( .A1(\DP_OP_487J11_125_9213/n18 ), .A2(
        \DP_OP_487J11_125_9213/n47 ), .Z(N1466) );
  XOR2D1BWP U8691 ( .A1(\DP_OP_487J11_125_9213/n17 ), .A2(
        \DP_OP_487J11_125_9213/n46 ), .Z(N1467) );
  OAI211D1BWP U8692 ( .A1(N1483), .A2(N1457), .B(N1469), .C(N1468), .ZN(n4136)
         );
  XOR2D1BWP U8693 ( .A1(\DP_OP_487J11_125_9213/n16 ), .A2(
        \DP_OP_487J11_125_9213/n45 ), .Z(N1468) );
  XOR2D1BWP U8694 ( .A1(\DP_OP_487J11_125_9213/n15 ), .A2(
        \DP_OP_487J11_125_9213/n44 ), .Z(N1469) );
  XOR2D1BWP U8695 ( .A1(\DP_OP_487J11_125_9213/n56 ), .A2(\C1/Z_0 ), .Z(N1457)
         );
  OAI211D1BWP U8696 ( .A1(N1470), .A2(n4374), .B(N1461), .C(N1459), .ZN(n4137)
         );
  XOR2D1BWP U8697 ( .A1(\DP_OP_487J11_125_9213/n25 ), .A2(
        \DP_OP_487J11_125_9213/n54 ), .Z(N1459) );
  XOR2D1BWP U8698 ( .A1(\DP_OP_487J11_125_9213/n23 ), .A2(
        \DP_OP_487J11_125_9213/n52 ), .Z(N1461) );
  AOI22D1BWP U8699 ( .A1(N1483), .A2(N1471), .B1(N1470), .B2(n4341), .ZN(n4139) );
  AOI21D1BWP U8700 ( .A1(n4151), .A2(n4636), .B(n4150), .ZN(n4354) );
  OAI31D1BWP U8701 ( .A1(n4359), .A2(n4149), .A3(n4148), .B(n4147), .ZN(n4150)
         );
  AOI22D1BWP U8702 ( .A1(N1483), .A2(N1476), .B1(N1475), .B2(n4341), .ZN(n4147) );
  NR2XD0BWP U8703 ( .A1(n4866), .A2(n4376), .ZN(n4373) );
  MUX2ND0BWP U8704 ( .I0(N1470), .I1(N1471), .S(n4355), .ZN(n4149) );
  XOR2D1BWP U8705 ( .A1(\DP_OP_487J11_125_9213/n13 ), .A2(
        \DP_OP_487J11_125_9213/n42 ), .Z(N1471) );
  NR2XD0BWP U8706 ( .A1(n4369), .A2(n4637), .ZN(n4636) );
  MUX2ND0BWP U8707 ( .I0(n4339), .I1(n4140), .S(n4359), .ZN(n4151) );
  MUX2ND0BWP U8708 ( .I0(N1472), .I1(N1473), .S(n4355), .ZN(n4140) );
  MUX2ND0BWP U8709 ( .I0(N1474), .I1(N1475), .S(n4355), .ZN(n4339) );
  AOI21D1BWP U8710 ( .A1(n4366), .A2(n4365), .B(n4364), .ZN(n4891) );
  MUX2ND0BWP U8711 ( .I0(n4363), .I1(n4362), .S(n4361), .ZN(n4364) );
  NR2XD0BWP U8712 ( .A1(n4374), .A2(n4360), .ZN(n4361) );
  XNR3D1BWP U8713 ( .A1(n4359), .A2(n4362), .A3(n4358), .ZN(n4365) );
  NR2XD0BWP U8714 ( .A1(N1481), .A2(n4101), .ZN(n4355) );
  MUX2ND0BWP U8715 ( .I0(result[10]), .I1(scalarToLoad[10]), .S(\intadd_34/n1 ), .ZN(n4360) );
  MUX2ND0BWP U8716 ( .I0(result[11]), .I1(scalarToLoad[11]), .S(\intadd_34/CO ), .ZN(n4120) );
  NR2XD0BWP U8717 ( .A1(N1481), .A2(n4143), .ZN(n4359) );
  ND3D1BWP U8718 ( .A1(n4097), .A2(n4146), .A3(n4374), .ZN(n4337) );
  NR2XD0BWP U8719 ( .A1(n4095), .A2(N1481), .ZN(n4090) );
  OR2XD1BWP U8720 ( .A1(N1480), .A2(N1479), .Z(n4095) );
  NR2XD0BWP U8721 ( .A1(N1476), .A2(N1475), .ZN(n4094) );
  NR2XD0BWP U8722 ( .A1(N1478), .A2(N1477), .ZN(n4096) );
  NR2XD0BWP U8723 ( .A1(n4093), .A2(N1472), .ZN(n4097) );
  OAI22D1BWP U8724 ( .A1(\intadd_34/CO ), .A2(n4231), .B1(n4230), .B2(n3676), 
        .ZN(\C3/Z_14 ) );
  AOI22D1BWP U8725 ( .A1(n4246), .A2(n4289), .B1(n4302), .B2(n4288), .ZN(n4230) );
  AOI222D1BWP U8726 ( .A1(n4311), .A2(n4242), .B1(n4285), .B2(n4273), .C1(
        n4286), .C2(n4302), .ZN(n4231) );
  OAI22D1BWP U8727 ( .A1(\intadd_34/CO ), .A2(n4239), .B1(n4238), .B2(n3676), 
        .ZN(\C3/Z_13 ) );
  AOI22D1BWP U8728 ( .A1(n4246), .A2(n4295), .B1(n4320), .B2(n4294), .ZN(n4238) );
  AOI22D1BWP U8729 ( .A1(n4246), .A2(n4293), .B1(n4320), .B2(n4292), .ZN(n4239) );
  OAI22D1BWP U8730 ( .A1(\intadd_34/n1 ), .A2(n4244), .B1(n4243), .B2(n3676), 
        .ZN(\C3/Z_12 ) );
  AOI222D1BWP U8731 ( .A1(n4242), .A2(n4332), .B1(n4273), .B2(n4301), .C1(
        n4320), .C2(n4300), .ZN(n4243) );
  AOI222D1BWP U8732 ( .A1(n4299), .A2(n4273), .B1(n4242), .B2(n4330), .C1(
        n4298), .C2(n4320), .ZN(n4244) );
  OAI22D1BWP U8733 ( .A1(\intadd_34/CO ), .A2(n4248), .B1(n4247), .B2(n3676), 
        .ZN(\C3/Z_11 ) );
  AOI22D1BWP U8734 ( .A1(n4246), .A2(n4308), .B1(n4320), .B2(n4307), .ZN(n4247) );
  AOI22D1BWP U8735 ( .A1(n4273), .A2(n4306), .B1(n4320), .B2(n4305), .ZN(n4248) );
  OAI22D1BWP U8736 ( .A1(\intadd_34/CO ), .A2(n4251), .B1(n4250), .B2(n3676), 
        .ZN(\C3/Z_10 ) );
  AOI22D1BWP U8737 ( .A1(n4273), .A2(n4313), .B1(n4320), .B2(n4314), .ZN(n4250) );
  AOI22D1BWP U8738 ( .A1(n4320), .A2(n4312), .B1(n4273), .B2(n4311), .ZN(n4251) );
  OAI22D1BWP U8739 ( .A1(\intadd_34/CO ), .A2(n4265), .B1(n4264), .B2(n3676), 
        .ZN(\C3/Z_9 ) );
  AOI21D1BWP U8740 ( .A1(n4315), .A2(n4326), .B(n4263), .ZN(n4264) );
  OAI22D1BWP U8741 ( .A1(n4324), .A2(n4272), .B1(n4262), .B2(n4321), .ZN(n4263) );
  OA222D1BWP U8742 ( .A1(n4260), .A2(n4259), .B1(n4323), .B2(n4258), .C1(n4257), .C2(n4256), .Z(n4265) );
  AOI21D1BWP U8743 ( .A1(n4320), .A2(n4255), .B(n4333), .ZN(n4256) );
  OAI22D1BWP U8744 ( .A1(\intadd_34/CO ), .A2(n4278), .B1(n4277), .B2(n3676), 
        .ZN(\C3/Z_8 ) );
  AOI222D1BWP U8745 ( .A1(n4276), .A2(n4275), .B1(n4315), .B2(n4274), .C1(
        n4273), .C2(n4332), .ZN(n4277) );
  OAI21D1BWP U8746 ( .A1(n4272), .A2(n4271), .B(n4322), .ZN(n4276) );
  AOI222D1BWP U8747 ( .A1(n4270), .A2(n4269), .B1(n4287), .B2(n4268), .C1(
        n4273), .C2(n4330), .ZN(n4278) );
  OAI21D1BWP U8748 ( .A1(n4266), .A2(n4272), .B(n4322), .ZN(n4270) );
  OAI22D1BWP U8749 ( .A1(\intadd_34/CO ), .A2(n4284), .B1(n4283), .B2(n3676), 
        .ZN(\C3/Z_7 ) );
  AOI22D1BWP U8750 ( .A1(n4320), .A2(n4282), .B1(n4287), .B2(n4281), .ZN(n4283) );
  AOI222D1BWP U8751 ( .A1(n4306), .A2(n4302), .B1(n4280), .B2(n4333), .C1(
        n4279), .C2(n4287), .ZN(n4284) );
  OAI22D1BWP U8752 ( .A1(\intadd_34/CO ), .A2(n4291), .B1(n4290), .B2(n3676), 
        .ZN(\C3/Z_6 ) );
  AOI22D1BWP U8753 ( .A1(n4320), .A2(n4289), .B1(n4288), .B2(n4287), .ZN(n4290) );
  MUX2ND0BWP U8754 ( .I0(n4249), .I1(n4229), .S(\intadd_34/SUM[1] ), .ZN(n4289) );
  AOI222D1BWP U8755 ( .A1(n4311), .A2(n4302), .B1(n4286), .B2(n4287), .C1(
        n4333), .C2(n4285), .ZN(n4291) );
  NR2XD0BWP U8756 ( .A1(n4323), .A2(\intadd_34/SUM[1] ), .ZN(n4287) );
  OAI22D1BWP U8757 ( .A1(\intadd_34/CO ), .A2(n4297), .B1(n4296), .B2(n3676), 
        .ZN(\C3/Z_5 ) );
  AOI22D1BWP U8758 ( .A1(n4320), .A2(n4295), .B1(n4315), .B2(n4294), .ZN(n4296) );
  AOI211XD0BWP U8759 ( .A1(n4710), .A2(n4237), .B(n4236), .C(n4235), .ZN(n4295) );
  OAI31D1BWP U8760 ( .A1(n4711), .A2(n4254), .A3(n4237), .B(n4234), .ZN(n4235)
         );
  NR2XD0BWP U8761 ( .A1(n4261), .A2(\intadd_34/SUM[1] ), .ZN(n4236) );
  AOI22D1BWP U8762 ( .A1(n4320), .A2(n4293), .B1(n4315), .B2(n4292), .ZN(n4297) );
  MUX2ND0BWP U8763 ( .I0(n4252), .I1(n4233), .S(\intadd_34/SUM[1] ), .ZN(n4293) );
  OAI22D1BWP U8764 ( .A1(\intadd_34/CO ), .A2(n4304), .B1(n4303), .B2(n3676), 
        .ZN(\C3/Z_4 ) );
  AOI222D1BWP U8765 ( .A1(n4302), .A2(n4332), .B1(n4333), .B2(n4301), .C1(
        n4315), .C2(n4300), .ZN(n4303) );
  AOI222D1BWP U8766 ( .A1(n4299), .A2(n4333), .B1(n4302), .B2(n4330), .C1(
        n4298), .C2(n4315), .ZN(n4304) );
  OAI22D1BWP U8767 ( .A1(\intadd_34/CO ), .A2(n4310), .B1(n4309), .B2(n3676), 
        .ZN(\C3/Z_3 ) );
  AOI22D1BWP U8768 ( .A1(n4320), .A2(n4308), .B1(n4315), .B2(n4307), .ZN(n4309) );
  NR2XD0BWP U8769 ( .A1(n4245), .A2(n4254), .ZN(n4308) );
  AOI22D1BWP U8770 ( .A1(n4333), .A2(n4306), .B1(n4315), .B2(n4305), .ZN(n4310) );
  OAI22D1BWP U8771 ( .A1(\intadd_34/CO ), .A2(n4317), .B1(n4316), .B2(n3676), 
        .ZN(\C3/Z_2 ) );
  AOI22D1BWP U8772 ( .A1(n4315), .A2(n4314), .B1(n4333), .B2(n4313), .ZN(n4316) );
  AOI22D1BWP U8773 ( .A1(n4315), .A2(n4312), .B1(n4333), .B2(n4311), .ZN(n4317) );
  AO222D1BWP U8774 ( .A1(scalarToLoad[1]), .A2(n4227), .B1(scalarToLoad[2]), 
        .B2(n4226), .C1(scalarToLoad[0]), .C2(n4228), .Z(n4311) );
  OAI22D1BWP U8775 ( .A1(\intadd_34/n1 ), .A2(n4328), .B1(n4327), .B2(n3676), 
        .ZN(\C3/Z_1 ) );
  AOI31D1BWP U8776 ( .A1(\intadd_34/SUM[2] ), .A2(\intadd_34/SUM[3] ), .A3(
        n4326), .B(n4325), .ZN(n4327) );
  OAI22D1BWP U8777 ( .A1(n4324), .A2(n4323), .B1(n4322), .B2(n4321), .ZN(n4325) );
  AOI22D1BWP U8778 ( .A1(n4320), .A2(n4319), .B1(\intadd_34/SUM[3] ), .B2(
        n4318), .ZN(n4328) );
  NR2XD0BWP U8779 ( .A1(n4252), .A2(n4254), .ZN(n4319) );
  OAI211D1BWP U8780 ( .A1(scalarToLoad[1]), .A2(n4638), .B(\intadd_34/SUM[0] ), 
        .C(n4232), .ZN(n4252) );
  OAI22D1BWP U8781 ( .A1(\intadd_34/n1 ), .A2(n4335), .B1(n4334), .B2(n3676), 
        .ZN(\C3/Z_0 ) );
  AOI22D1BWP U8782 ( .A1(n4333), .A2(n4332), .B1(\intadd_34/SUM[3] ), .B2(
        n4331), .ZN(n4334) );
  NR2XD0BWP U8783 ( .A1(n4241), .A2(n6004), .ZN(n4332) );
  AOI22D1BWP U8784 ( .A1(n4333), .A2(n4330), .B1(\intadd_34/SUM[3] ), .B2(
        n4329), .ZN(n4335) );
  NR2XD0BWP U8785 ( .A1(n4240), .A2(n4241), .ZN(n4330) );
  NR2XD0BWP U8786 ( .A1(n4272), .A2(n4254), .ZN(n4333) );
  MUX2ND0BWP U8787 ( .I0(n4245), .I1(n4224), .S(\intadd_34/SUM[1] ), .ZN(n4282) );
  MUX2D1BWP U8788 ( .I0(n4709), .I1(n4710), .S(\intadd_34/SUM[0] ), .Z(n4245)
         );
  AOI22D1BWP U8789 ( .A1(n4638), .A2(result[0]), .B1(result[1]), .B2(n4706), 
        .ZN(n4709) );
  NR2XD0BWP U8790 ( .A1(n4272), .A2(\intadd_34/SUM[1] ), .ZN(n4302) );
  NR2XD0BWP U8791 ( .A1(n4254), .A2(n4260), .ZN(n4273) );
  AOI22D1BWP U8792 ( .A1(scalarToLoad[1]), .A2(n4228), .B1(scalarToLoad[0]), 
        .B2(n4219), .ZN(n4220) );
  AOI22D1BWP U8793 ( .A1(n4227), .A2(scalarToLoad[2]), .B1(n4226), .B2(
        scalarToLoad[3]), .ZN(n4221) );
  OAI22D1BWP U8794 ( .A1(\intadd_34/n1 ), .A2(n4643), .B1(n4162), .B2(n3676), 
        .ZN(\C2/Z_16 ) );
  OAI31D1BWP U8795 ( .A1(\intadd_34/SUM[3] ), .A2(n3676), .A3(n4218), .B(n4217), .ZN(\C3/Z_16 ) );
  OA211D1BWP U8796 ( .A1(n4299), .A2(n4215), .B(n4214), .C(n4269), .Z(n4329)
         );
  OAI21D1BWP U8797 ( .A1(\intadd_34/SUM[1] ), .A2(n4267), .B(
        \intadd_34/SUM[2] ), .ZN(n4214) );
  AOI22D1BWP U8798 ( .A1(scalarToLoad[1]), .A2(n4219), .B1(scalarToLoad[2]), 
        .B2(n4228), .ZN(n4211) );
  AOI22D1BWP U8799 ( .A1(n4227), .A2(scalarToLoad[3]), .B1(n4226), .B2(
        scalarToLoad[4]), .ZN(n4212) );
  AOI21D1BWP U8800 ( .A1(n4210), .A2(n4271), .B(n4209), .ZN(n4331) );
  AOI21D1BWP U8801 ( .A1(n4253), .A2(n4275), .B(n4274), .ZN(n4209) );
  MUX2ND0BWP U8802 ( .I0(n4705), .I1(n4208), .S(\intadd_34/SUM[0] ), .ZN(n4301) );
  OAI22D1BWP U8803 ( .A1(n4706), .A2(result[1]), .B1(result[2]), .B2(n4638), 
        .ZN(n4705) );
  OAI22D1BWP U8804 ( .A1(\intadd_34/CO ), .A2(n4668), .B1(n4158), .B2(n3676), 
        .ZN(\C2/Z_17 ) );
  NR2XD0BWP U8805 ( .A1(\intadd_34/CO ), .A2(\intadd_34/SUM[3] ), .ZN(n4216)
         );
  AOI211XD0BWP U8806 ( .A1(\intadd_34/SUM[2] ), .A2(n4258), .B(n4206), .C(
        n4257), .ZN(n4318) );
  NR2XD0BWP U8807 ( .A1(n4205), .A2(n4254), .ZN(n4257) );
  NR2XD0BWP U8808 ( .A1(n4215), .A2(n4255), .ZN(n4206) );
  NR2XD0BWP U8809 ( .A1(n4204), .A2(n4203), .ZN(n4255) );
  OAI22D1BWP U8810 ( .A1(scalarToLoad[5]), .A2(n4241), .B1(scalarToLoad[4]), 
        .B2(n4202), .ZN(n4203) );
  OAI22D1BWP U8811 ( .A1(scalarToLoad[2]), .A2(n4201), .B1(scalarToLoad[3]), 
        .B2(n4200), .ZN(n4204) );
  AOI21D1BWP U8812 ( .A1(\intadd_34/SUM[1] ), .A2(n4199), .B(n4198), .ZN(n4324) );
  OAI22D1BWP U8813 ( .A1(n4710), .A2(n4234), .B1(n4237), .B2(n4197), .ZN(n4198) );
  OAI22D1BWP U8814 ( .A1(n4706), .A2(result[2]), .B1(result[3]), .B2(n4638), 
        .ZN(n4710) );
  MUX2ND0BWP U8815 ( .I0(n4196), .I1(n4708), .S(\intadd_34/SUM[0] ), .ZN(n4199) );
  OAI22D1BWP U8816 ( .A1(\intadd_34/n1 ), .A2(n6011), .B1(n4157), .B2(n3676), 
        .ZN(\C2/Z_18 ) );
  AO22D1BWP U8817 ( .A1(n4194), .A2(n4314), .B1(n4193), .B2(n4312), .Z(
        \C3/Z_18 ) );
  MUX2ND0BWP U8818 ( .I0(n4192), .I1(n4191), .S(\intadd_34/SUM[1] ), .ZN(n4312) );
  NR2XD0BWP U8819 ( .A1(n4190), .A2(n4189), .ZN(n4285) );
  OAI22D1BWP U8820 ( .A1(scalarToLoad[5]), .A2(n4202), .B1(scalarToLoad[6]), 
        .B2(n4241), .ZN(n4189) );
  OAI22D1BWP U8821 ( .A1(scalarToLoad[4]), .A2(n4200), .B1(scalarToLoad[3]), 
        .B2(n4201), .ZN(n4190) );
  MUX2ND0BWP U8822 ( .I0(n4229), .I1(n4188), .S(\intadd_34/SUM[1] ), .ZN(n4314) );
  MUX2ND0BWP U8823 ( .I0(n4703), .I1(n4704), .S(\intadd_34/SUM[0] ), .ZN(n4229) );
  AOI22D1BWP U8824 ( .A1(n4638), .A2(n6011), .B1(n4665), .B2(n4706), .ZN(n4703) );
  OAI22D1BWP U8825 ( .A1(\intadd_34/CO ), .A2(n4665), .B1(n4154), .B2(n3676), 
        .ZN(\C2/Z_19 ) );
  AO22D1BWP U8826 ( .A1(n4305), .A2(n4193), .B1(n4307), .B2(n4194), .Z(
        \C3/Z_19 ) );
  MUX2ND0BWP U8827 ( .I0(n4224), .I1(n4225), .S(\intadd_34/SUM[1] ), .ZN(n4307) );
  MUX2ND0BWP U8828 ( .I0(n4711), .I1(n4707), .S(\intadd_34/SUM[0] ), .ZN(n4224) );
  AOI22D1BWP U8829 ( .A1(n4638), .A2(n4665), .B1(n4664), .B2(n4706), .ZN(n4711) );
  MUX2ND0BWP U8830 ( .I0(n4222), .I1(n4223), .S(\intadd_34/SUM[1] ), .ZN(n4305) );
  OA211D1BWP U8831 ( .A1(n4241), .A2(n4187), .B(n4186), .C(n4185), .Z(n4222)
         );
  AOI22D1BWP U8832 ( .A1(n4228), .A2(scalarToLoad[5]), .B1(n4219), .B2(
        scalarToLoad[4]), .ZN(n4186) );
  MUX2ND0BWP U8833 ( .I0(n4213), .I1(n4267), .S(\intadd_34/SUM[1] ), .ZN(n4298) );
  AO211D1BWP U8834 ( .A1(n4227), .A2(n4187), .B(n4184), .C(n4183), .Z(n4213)
         );
  OAI22D1BWP U8835 ( .A1(scalarToLoad[5]), .A2(n4201), .B1(scalarToLoad[6]), 
        .B2(n4200), .ZN(n4183) );
  NR2XD0BWP U8836 ( .A1(n4241), .A2(scalarToLoad[8]), .ZN(n4184) );
  AOI22D1BWP U8837 ( .A1(n4638), .A2(n4664), .B1(n4661), .B2(n4706), .ZN(n4704) );
  OAI22D1BWP U8838 ( .A1(n4661), .A2(\intadd_34/CO ), .B1(n4133), .B2(n3676), 
        .ZN(\C2/Z_21 ) );
  AO22D1BWP U8839 ( .A1(n4193), .A2(n4292), .B1(n4194), .B2(n4294), .Z(
        \C3/Z_21 ) );
  AOI222D1BWP U8840 ( .A1(n4181), .A2(\intadd_34/SUM[1] ), .B1(
        \intadd_34/SUM[0] ), .B2(n4708), .C1(n4196), .C2(n4180), .ZN(n4294) );
  AOI22D1BWP U8841 ( .A1(n4638), .A2(n4661), .B1(n4655), .B2(n4706), .ZN(n4707) );
  MUX2D1BWP U8842 ( .I0(n4205), .I1(n4179), .S(\intadd_34/SUM[1] ), .Z(n4292)
         );
  AOI22D1BWP U8843 ( .A1(scalarToLoad[7]), .A2(n4228), .B1(n4219), .B2(
        scalarToLoad[6]), .ZN(n4177) );
  AOI22D1BWP U8844 ( .A1(n4227), .A2(scalarToLoad[8]), .B1(n4226), .B2(
        scalarToLoad[9]), .ZN(n4178) );
  NR2XD0BWP U8845 ( .A1(n4237), .A2(n4638), .ZN(n4226) );
  OAI22D1BWP U8846 ( .A1(n4655), .A2(\intadd_34/CO ), .B1(n3676), .B2(n4187), 
        .ZN(\C2/Z_22 ) );
  OAI22D1BWP U8847 ( .A1(n4191), .A2(n4176), .B1(n4188), .B2(n4175), .ZN(
        \C3/Z_22 ) );
  AOI21D1BWP U8848 ( .A1(\intadd_34/SUM[0] ), .A2(n4174), .B(n4173), .ZN(n4288) );
  OAI22D1BWP U8849 ( .A1(\intadd_34/SUM[0] ), .A2(n4702), .B1(result[9]), .B2(
        n4202), .ZN(n4173) );
  AOI22D1BWP U8850 ( .A1(n4638), .A2(n4655), .B1(n4652), .B2(n4706), .ZN(n4702) );
  AOI211XD0BWP U8851 ( .A1(n4219), .A2(n4187), .B(n4172), .C(n4171), .ZN(n4286) );
  OAI22D1BWP U8852 ( .A1(scalarToLoad[9]), .A2(n4202), .B1(scalarToLoad[8]), 
        .B2(n4200), .ZN(n4171) );
  NR3D0BWP U8853 ( .A1(n4699), .A2(n4237), .A3(n4170), .ZN(n4172) );
  OAI22D1BWP U8854 ( .A1(n4652), .A2(\intadd_34/CO ), .B1(n4106), .B2(n3676), 
        .ZN(\C2/Z_23 ) );
  OAI22D1BWP U8855 ( .A1(n4225), .A2(n4175), .B1(n4223), .B2(n4176), .ZN(
        \C3/Z_23 ) );
  AOI222D1BWP U8856 ( .A1(n4170), .A2(n4227), .B1(n4219), .B2(scalarToLoad[8]), 
        .C1(n4228), .C2(scalarToLoad[9]), .ZN(n4223) );
  NR2XD0BWP U8857 ( .A1(n4638), .A2(\intadd_34/SUM[0] ), .ZN(n4228) );
  OAI22D1BWP U8858 ( .A1(n4706), .A2(result[8]), .B1(result[9]), .B2(n4638), 
        .ZN(n4708) );
  NR2XD0BWP U8859 ( .A1(n4237), .A2(n4706), .ZN(n4227) );
  OAI22D1BWP U8860 ( .A1(n4651), .A2(\intadd_34/n1 ), .B1(n4088), .B2(n3676), 
        .ZN(\C2/Z_24 ) );
  AOI211XD0BWP U8861 ( .A1(n4638), .A2(n4651), .B(\intadd_34/SUM[0] ), .C(
        n4174), .ZN(n4182) );
  NR2XD0BWP U8862 ( .A1(n4169), .A2(n3615), .ZN(n4174) );
  NR2XD0BWP U8863 ( .A1(n4260), .A2(\intadd_34/SUM[1] ), .ZN(n4242) );
  OAI211D1BWP U8864 ( .A1(scalarToLoad[9]), .A2(n4706), .B(n4237), .C(n4168), 
        .ZN(n4267) );
  OAI22D1BWP U8865 ( .A1(\intadd_34/CO ), .A2(n4087), .B1(n4167), .B2(n3676), 
        .ZN(\C2/Z_25 ) );
  NR2XD0BWP U8866 ( .A1(n4260), .A2(n3676), .ZN(n4194) );
  NR2XD0BWP U8867 ( .A1(n4181), .A2(\intadd_34/SUM[1] ), .ZN(n4326) );
  NR4D0BWP U8868 ( .A1(result[10]), .A2(result[12]), .A3(result[11]), .A4(
        result[13]), .ZN(n4085) );
  NR2XD0BWP U8869 ( .A1(n4260), .A2(\intadd_34/CO ), .ZN(n4193) );
  FA1D0BWP U8870 ( .A(\intadd_34/A[1] ), .B(scalarToLoad[12]), .CI(
        \intadd_34/n4 ), .CO(\intadd_34/n3 ), .S(\intadd_34/SUM[1] ) );
  NR2XD0BWP U8871 ( .A1(n4201), .A2(n4167), .ZN(n4179) );
  ND4D1BWP U8872 ( .A1(n4086), .A2(n3615), .A3(n3638), .A4(n3655), .ZN(n4170)
         );
  NR2XD0BWP U8873 ( .A1(scalarToLoad[12]), .A2(scalarToLoad[11]), .ZN(n4086)
         );
  FA1D0BWP U8874 ( .A(\intadd_34/A[0] ), .B(scalarToLoad[11]), .CI(
        \intadd_34/CI ), .CO(\intadd_34/n4 ), .S(\intadd_34/SUM[0] ) );
  OA21D1BWP U8875 ( .A1(result[10]), .A2(n3615), .B(\intadd_34/CI ), .Z(n4638)
         );
  OAI211D1BWP U8876 ( .A1(n6038), .A2(n4643), .B(n6006), .C(n6005), .ZN(
        \srf/N38 ) );
  AOI22D1BWP U8877 ( .A1(n4065), .A2(Addr[1]), .B1(n6034), .B2(\srf/N34 ), 
        .ZN(n6006) );
  ND4D1BWP U8878 ( .A1(n8142), .A2(n8143), .A3(n8144), .A4(n8145), .ZN(
        \srf/N34 ) );
  AOI22D1BWP U8879 ( .A1(n8136), .A2(\srf/regTable[5][1] ), .B1(n8137), .B2(
        \srf/regTable[7][1] ), .ZN(n8145) );
  AOI22D1BWP U8880 ( .A1(n8134), .A2(\srf/regTable[4][1] ), .B1(n8135), .B2(
        \srf/regTable[6][1] ), .ZN(n8144) );
  AOI22D1BWP U8881 ( .A1(n8131), .A2(\srf/regTable[1][1] ), .B1(n8133), .B2(
        \srf/regTable[3][1] ), .ZN(n8143) );
  AOI22D1BWP U8882 ( .A1(n8127), .A2(\srf/regTable[0][1] ), .B1(n8129), .B2(
        \srf/regTable[2][1] ), .ZN(n8142) );
  OAI211D1BWP U8883 ( .A1(n6038), .A2(n6004), .B(n6003), .C(n6002), .ZN(
        \srf/N37 ) );
  AOI22D1BWP U8884 ( .A1(n4065), .A2(Addr[0]), .B1(n6034), .B2(\srf/N35 ), 
        .ZN(n6003) );
  ND4D1BWP U8885 ( .A1(n8138), .A2(n8139), .A3(n8140), .A4(n8141), .ZN(
        \srf/N35 ) );
  AOI22D1BWP U8886 ( .A1(n8136), .A2(\srf/regTable[5][0] ), .B1(n8137), .B2(
        \srf/regTable[7][0] ), .ZN(n8141) );
  AOI22D1BWP U8887 ( .A1(n8134), .A2(\srf/regTable[4][0] ), .B1(n8135), .B2(
        \srf/regTable[6][0] ), .ZN(n8140) );
  AOI22D1BWP U8888 ( .A1(n8131), .A2(\srf/regTable[1][0] ), .B1(n8133), .B2(
        \srf/regTable[3][0] ), .ZN(n8139) );
  AOI22D1BWP U8889 ( .A1(n8127), .A2(\srf/regTable[0][0] ), .B1(n8129), .B2(
        \srf/regTable[2][0] ), .ZN(n8138) );
  OAI211D1BWP U8890 ( .A1(n6038), .A2(n6037), .B(n6036), .C(n6035), .ZN(
        \srf/N52 ) );
  AOI22D1BWP U8891 ( .A1(n4065), .A2(Addr[15]), .B1(n6034), .B2(\srf/N20 ), 
        .ZN(n6036) );
  ND4D1BWP U8892 ( .A1(n8198), .A2(n8199), .A3(n8200), .A4(n8201), .ZN(
        \srf/N20 ) );
  AOI22D1BWP U8893 ( .A1(n8136), .A2(\srf/regTable[5][15] ), .B1(n8137), .B2(
        \srf/regTable[7][15] ), .ZN(n8201) );
  AOI22D1BWP U8894 ( .A1(n8134), .A2(\srf/regTable[4][15] ), .B1(n8135), .B2(
        \srf/regTable[6][15] ), .ZN(n8200) );
  AOI22D1BWP U8895 ( .A1(n8131), .A2(\srf/regTable[1][15] ), .B1(n8133), .B2(
        \srf/regTable[3][15] ), .ZN(n8199) );
  AOI22D1BWP U8896 ( .A1(n8127), .A2(\srf/regTable[0][15] ), .B1(n8129), .B2(
        \srf/regTable[2][15] ), .ZN(n8198) );
  OAI211D1BWP U8897 ( .A1(n6038), .A2(\intadd_34/A[3] ), .B(n6033), .C(n6032), 
        .ZN(\srf/N51 ) );
  AOI22D1BWP U8898 ( .A1(n4065), .A2(Addr[14]), .B1(n6034), .B2(\srf/N21 ), 
        .ZN(n6033) );
  ND4D1BWP U8899 ( .A1(n8194), .A2(n8195), .A3(n8196), .A4(n8197), .ZN(
        \srf/N21 ) );
  AOI22D1BWP U8900 ( .A1(n8136), .A2(\srf/regTable[5][14] ), .B1(n8137), .B2(
        \srf/regTable[7][14] ), .ZN(n8197) );
  AOI22D1BWP U8901 ( .A1(n8134), .A2(\srf/regTable[4][14] ), .B1(n8135), .B2(
        \srf/regTable[6][14] ), .ZN(n8196) );
  AOI22D1BWP U8902 ( .A1(n8131), .A2(\srf/regTable[1][14] ), .B1(n8133), .B2(
        \srf/regTable[3][14] ), .ZN(n8195) );
  AOI22D1BWP U8903 ( .A1(n8127), .A2(\srf/regTable[0][14] ), .B1(n8129), .B2(
        \srf/regTable[2][14] ), .ZN(n8194) );
  INVD1BWP U8904 ( .I(result[14]), .ZN(\intadd_34/A[3] ) );
  OAI211D1BWP U8905 ( .A1(n6038), .A2(\intadd_34/A[2] ), .B(n6031), .C(n6030), 
        .ZN(\srf/N50 ) );
  AOI22D1BWP U8906 ( .A1(n4065), .A2(Addr[13]), .B1(n6034), .B2(\srf/N22 ), 
        .ZN(n6031) );
  ND4D1BWP U8907 ( .A1(n8190), .A2(n8191), .A3(n8192), .A4(n8193), .ZN(
        \srf/N22 ) );
  AOI22D1BWP U8908 ( .A1(n8136), .A2(\srf/regTable[5][13] ), .B1(n8137), .B2(
        \srf/regTable[7][13] ), .ZN(n8193) );
  AOI22D1BWP U8909 ( .A1(n8134), .A2(\srf/regTable[4][13] ), .B1(n8135), .B2(
        \srf/regTable[6][13] ), .ZN(n8192) );
  AOI22D1BWP U8910 ( .A1(n8131), .A2(\srf/regTable[1][13] ), .B1(n8133), .B2(
        \srf/regTable[3][13] ), .ZN(n8191) );
  AOI22D1BWP U8911 ( .A1(n8127), .A2(\srf/regTable[0][13] ), .B1(n8129), .B2(
        \srf/regTable[2][13] ), .ZN(n8190) );
  OAI211D1BWP U8912 ( .A1(n6038), .A2(\intadd_34/A[1] ), .B(n6029), .C(n6028), 
        .ZN(\srf/N49 ) );
  AOI22D1BWP U8913 ( .A1(n4065), .A2(Addr[12]), .B1(n6034), .B2(\srf/N23 ), 
        .ZN(n6029) );
  ND4D1BWP U8914 ( .A1(n8186), .A2(n8187), .A3(n8188), .A4(n8189), .ZN(
        \srf/N23 ) );
  AOI22D1BWP U8915 ( .A1(n8136), .A2(\srf/regTable[5][12] ), .B1(n8137), .B2(
        \srf/regTable[7][12] ), .ZN(n8189) );
  AOI22D1BWP U8916 ( .A1(n8134), .A2(\srf/regTable[4][12] ), .B1(n8135), .B2(
        \srf/regTable[6][12] ), .ZN(n8188) );
  AOI22D1BWP U8917 ( .A1(n8131), .A2(\srf/regTable[1][12] ), .B1(n8133), .B2(
        \srf/regTable[3][12] ), .ZN(n8187) );
  AOI22D1BWP U8918 ( .A1(n8127), .A2(\srf/regTable[0][12] ), .B1(n8129), .B2(
        \srf/regTable[2][12] ), .ZN(n8186) );
  OAI211D1BWP U8919 ( .A1(n6038), .A2(\intadd_34/A[0] ), .B(n6027), .C(n6026), 
        .ZN(\srf/N48 ) );
  AOI22D1BWP U8920 ( .A1(n4065), .A2(Addr[11]), .B1(n6034), .B2(\srf/N24 ), 
        .ZN(n6027) );
  ND4D1BWP U8921 ( .A1(n8182), .A2(n8183), .A3(n8184), .A4(n8185), .ZN(
        \srf/N24 ) );
  AOI22D1BWP U8922 ( .A1(n8136), .A2(\srf/regTable[5][11] ), .B1(n8137), .B2(
        \srf/regTable[7][11] ), .ZN(n8185) );
  AOI22D1BWP U8923 ( .A1(n8134), .A2(\srf/regTable[4][11] ), .B1(n8135), .B2(
        \srf/regTable[6][11] ), .ZN(n8184) );
  AOI22D1BWP U8924 ( .A1(n8131), .A2(\srf/regTable[1][11] ), .B1(n8133), .B2(
        \srf/regTable[3][11] ), .ZN(n8183) );
  AOI22D1BWP U8925 ( .A1(n8127), .A2(\srf/regTable[0][11] ), .B1(n8129), .B2(
        \srf/regTable[2][11] ), .ZN(n8182) );
  OAI211D1BWP U8926 ( .A1(n6038), .A2(n4699), .B(n6025), .C(n6024), .ZN(
        \srf/N47 ) );
  AOI22D1BWP U8927 ( .A1(n4065), .A2(Addr[10]), .B1(n6034), .B2(\srf/N25 ), 
        .ZN(n6025) );
  ND4D1BWP U8928 ( .A1(n8178), .A2(n8179), .A3(n8180), .A4(n8181), .ZN(
        \srf/N25 ) );
  AOI22D1BWP U8929 ( .A1(n8136), .A2(\srf/regTable[5][10] ), .B1(n8137), .B2(
        \srf/regTable[7][10] ), .ZN(n8181) );
  AOI22D1BWP U8930 ( .A1(n8134), .A2(\srf/regTable[4][10] ), .B1(n8135), .B2(
        \srf/regTable[6][10] ), .ZN(n8180) );
  AOI22D1BWP U8931 ( .A1(n8131), .A2(\srf/regTable[1][10] ), .B1(n8133), .B2(
        \srf/regTable[3][10] ), .ZN(n8179) );
  AOI22D1BWP U8932 ( .A1(n8127), .A2(\srf/regTable[0][10] ), .B1(n8129), .B2(
        \srf/regTable[2][10] ), .ZN(n8178) );
  OAI211D1BWP U8933 ( .A1(n6038), .A2(n4651), .B(n6023), .C(n6022), .ZN(
        \srf/N46 ) );
  AOI22D1BWP U8934 ( .A1(n4065), .A2(Addr[9]), .B1(n6034), .B2(\srf/N26 ), 
        .ZN(n6023) );
  ND4D1BWP U8935 ( .A1(n8174), .A2(n8175), .A3(n8176), .A4(n8177), .ZN(
        \srf/N26 ) );
  AOI22D1BWP U8936 ( .A1(n8136), .A2(\srf/regTable[5][9] ), .B1(n8137), .B2(
        \srf/regTable[7][9] ), .ZN(n8177) );
  AOI22D1BWP U8937 ( .A1(n8134), .A2(\srf/regTable[4][9] ), .B1(n8135), .B2(
        \srf/regTable[6][9] ), .ZN(n8176) );
  AOI22D1BWP U8938 ( .A1(n8131), .A2(\srf/regTable[1][9] ), .B1(n8133), .B2(
        \srf/regTable[3][9] ), .ZN(n8175) );
  AOI22D1BWP U8939 ( .A1(n8127), .A2(\srf/regTable[0][9] ), .B1(n8129), .B2(
        \srf/regTable[2][9] ), .ZN(n8174) );
  OAI211D1BWP U8940 ( .A1(n6038), .A2(n4652), .B(n6021), .C(n6020), .ZN(
        \srf/N45 ) );
  AOI22D1BWP U8941 ( .A1(n4065), .A2(Addr[8]), .B1(n6034), .B2(\srf/N27 ), 
        .ZN(n6021) );
  ND4D1BWP U8942 ( .A1(n8170), .A2(n8171), .A3(n8172), .A4(n8173), .ZN(
        \srf/N27 ) );
  AOI22D1BWP U8943 ( .A1(n8136), .A2(\srf/regTable[5][8] ), .B1(n8137), .B2(
        \srf/regTable[7][8] ), .ZN(n8173) );
  AOI22D1BWP U8944 ( .A1(n8134), .A2(\srf/regTable[4][8] ), .B1(n8135), .B2(
        \srf/regTable[6][8] ), .ZN(n8172) );
  AOI22D1BWP U8945 ( .A1(n8131), .A2(\srf/regTable[1][8] ), .B1(n8133), .B2(
        \srf/regTable[3][8] ), .ZN(n8171) );
  AOI22D1BWP U8946 ( .A1(n8127), .A2(\srf/regTable[0][8] ), .B1(n8129), .B2(
        \srf/regTable[2][8] ), .ZN(n8170) );
  OAI211D1BWP U8947 ( .A1(n6038), .A2(n4655), .B(n6019), .C(n6018), .ZN(
        \srf/N44 ) );
  AOI22D1BWP U8948 ( .A1(n4065), .A2(Addr[7]), .B1(n6034), .B2(\srf/N28 ), 
        .ZN(n6019) );
  ND4D1BWP U8949 ( .A1(n8166), .A2(n8167), .A3(n8168), .A4(n8169), .ZN(
        \srf/N28 ) );
  AOI22D1BWP U8950 ( .A1(n8136), .A2(\srf/regTable[5][7] ), .B1(n8137), .B2(
        \srf/regTable[7][7] ), .ZN(n8169) );
  AOI22D1BWP U8951 ( .A1(n8134), .A2(\srf/regTable[4][7] ), .B1(n8135), .B2(
        \srf/regTable[6][7] ), .ZN(n8168) );
  AOI22D1BWP U8952 ( .A1(n8131), .A2(\srf/regTable[1][7] ), .B1(n8133), .B2(
        \srf/regTable[3][7] ), .ZN(n8167) );
  AOI22D1BWP U8953 ( .A1(n8127), .A2(\srf/regTable[0][7] ), .B1(n8129), .B2(
        \srf/regTable[2][7] ), .ZN(n8166) );
  OAI211D1BWP U8954 ( .A1(n6038), .A2(n4661), .B(n6017), .C(n6016), .ZN(
        \srf/N43 ) );
  AOI22D1BWP U8955 ( .A1(n4065), .A2(Addr[6]), .B1(n6034), .B2(\srf/N29 ), 
        .ZN(n6017) );
  ND4D1BWP U8956 ( .A1(n8162), .A2(n8163), .A3(n8164), .A4(n8165), .ZN(
        \srf/N29 ) );
  AOI22D1BWP U8957 ( .A1(n8136), .A2(\srf/regTable[5][6] ), .B1(n8137), .B2(
        \srf/regTable[7][6] ), .ZN(n8165) );
  AOI22D1BWP U8958 ( .A1(n8134), .A2(\srf/regTable[4][6] ), .B1(n8135), .B2(
        \srf/regTable[6][6] ), .ZN(n8164) );
  AOI22D1BWP U8959 ( .A1(n8131), .A2(\srf/regTable[1][6] ), .B1(n8133), .B2(
        \srf/regTable[3][6] ), .ZN(n8163) );
  AOI22D1BWP U8960 ( .A1(n8127), .A2(\srf/regTable[0][6] ), .B1(n8129), .B2(
        \srf/regTable[2][6] ), .ZN(n8162) );
  OAI211D1BWP U8961 ( .A1(n6038), .A2(n4664), .B(n6015), .C(n6014), .ZN(
        \srf/N42 ) );
  AOI22D1BWP U8962 ( .A1(n4065), .A2(Addr[5]), .B1(n6034), .B2(\srf/N30 ), 
        .ZN(n6015) );
  ND4D1BWP U8963 ( .A1(n8158), .A2(n8159), .A3(n8160), .A4(n8161), .ZN(
        \srf/N30 ) );
  AOI22D1BWP U8964 ( .A1(n8136), .A2(\srf/regTable[5][5] ), .B1(n8137), .B2(
        \srf/regTable[7][5] ), .ZN(n8161) );
  AOI22D1BWP U8965 ( .A1(n8134), .A2(\srf/regTable[4][5] ), .B1(n8135), .B2(
        \srf/regTable[6][5] ), .ZN(n8160) );
  AOI22D1BWP U8966 ( .A1(n8131), .A2(\srf/regTable[1][5] ), .B1(n8133), .B2(
        \srf/regTable[3][5] ), .ZN(n8159) );
  AOI22D1BWP U8967 ( .A1(n8127), .A2(\srf/regTable[0][5] ), .B1(n8129), .B2(
        \srf/regTable[2][5] ), .ZN(n8158) );
  OAI211D1BWP U8968 ( .A1(n6038), .A2(n4665), .B(n6013), .C(n6012), .ZN(
        \srf/N41 ) );
  AOI22D1BWP U8969 ( .A1(n4065), .A2(Addr[4]), .B1(n6034), .B2(\srf/N31 ), 
        .ZN(n6013) );
  ND4D1BWP U8970 ( .A1(n8154), .A2(n8155), .A3(n8156), .A4(n8157), .ZN(
        \srf/N31 ) );
  AOI22D1BWP U8971 ( .A1(n8136), .A2(\srf/regTable[5][4] ), .B1(n8137), .B2(
        \srf/regTable[7][4] ), .ZN(n8157) );
  AOI22D1BWP U8972 ( .A1(n8134), .A2(\srf/regTable[4][4] ), .B1(n8135), .B2(
        \srf/regTable[6][4] ), .ZN(n8156) );
  AOI22D1BWP U8973 ( .A1(n8131), .A2(\srf/regTable[1][4] ), .B1(n8133), .B2(
        \srf/regTable[3][4] ), .ZN(n8155) );
  AOI22D1BWP U8974 ( .A1(n8127), .A2(\srf/regTable[0][4] ), .B1(n8129), .B2(
        \srf/regTable[2][4] ), .ZN(n8154) );
  OAI211D1BWP U8975 ( .A1(n6038), .A2(n6011), .B(n6010), .C(n6009), .ZN(
        \srf/N40 ) );
  AOI22D1BWP U8976 ( .A1(n4065), .A2(Addr[3]), .B1(n6034), .B2(\srf/N32 ), 
        .ZN(n6010) );
  ND4D1BWP U8977 ( .A1(n8150), .A2(n8151), .A3(n8152), .A4(n8153), .ZN(
        \srf/N32 ) );
  AOI22D1BWP U8978 ( .A1(n8136), .A2(\srf/regTable[5][3] ), .B1(n8137), .B2(
        \srf/regTable[7][3] ), .ZN(n8153) );
  AOI22D1BWP U8979 ( .A1(n8134), .A2(\srf/regTable[4][3] ), .B1(n8135), .B2(
        \srf/regTable[6][3] ), .ZN(n8152) );
  AOI22D1BWP U8980 ( .A1(n8131), .A2(\srf/regTable[1][3] ), .B1(n8133), .B2(
        \srf/regTable[3][3] ), .ZN(n8151) );
  AOI22D1BWP U8981 ( .A1(n8127), .A2(\srf/regTable[0][3] ), .B1(n8129), .B2(
        \srf/regTable[2][3] ), .ZN(n8150) );
  OAI211D1BWP U8982 ( .A1(n6038), .A2(n4668), .B(n6008), .C(n6007), .ZN(
        \srf/N39 ) );
  AOI22D1BWP U8983 ( .A1(n4065), .A2(Addr[2]), .B1(n6034), .B2(\srf/N33 ), 
        .ZN(n6008) );
  ND4D1BWP U8984 ( .A1(n8146), .A2(n8147), .A3(n8148), .A4(n8149), .ZN(
        \srf/N33 ) );
  AOI22D1BWP U8985 ( .A1(n8136), .A2(\srf/regTable[5][2] ), .B1(n8137), .B2(
        \srf/regTable[7][2] ), .ZN(n8149) );
  NR2XD0BWP U8986 ( .A1(n8132), .A2(n8202), .ZN(n8137) );
  NR2XD0BWP U8987 ( .A1(n8130), .A2(n8202), .ZN(n8136) );
  AOI22D1BWP U8988 ( .A1(n8134), .A2(\srf/regTable[4][2] ), .B1(n8135), .B2(
        \srf/regTable[6][2] ), .ZN(n8148) );
  NR2XD0BWP U8989 ( .A1(n8128), .A2(n8202), .ZN(n8135) );
  AOI22D1BWP U8990 ( .A1(n8131), .A2(\srf/regTable[1][2] ), .B1(n8133), .B2(
        \srf/regTable[3][2] ), .ZN(n8147) );
  NR2XD0BWP U8991 ( .A1(n8132), .A2(\srf/N17 ), .ZN(n8133) );
  NR2XD0BWP U8992 ( .A1(n8130), .A2(\srf/N17 ), .ZN(n8131) );
  AOI22D1BWP U8993 ( .A1(n8127), .A2(\srf/regTable[0][2] ), .B1(n8129), .B2(
        \srf/regTable[2][2] ), .ZN(n8146) );
  NR2XD0BWP U8994 ( .A1(n8128), .A2(\srf/N17 ), .ZN(n8129) );
  NR2XD0BWP U8995 ( .A1(n5247), .A2(n5248), .ZN(n5997) );
  AOI21D1BWP U8996 ( .A1(n4561), .A2(n6000), .B(n4468), .ZN(n5248) );
  ND3D1BWP U8997 ( .A1(n4572), .A2(n4661), .A3(n4057), .ZN(n4058) );
  NR3D0BWP U8998 ( .A1(n4988), .A2(n4642), .A3(n4074), .ZN(n4057) );
  ND4D1BWP U8999 ( .A1(result[10]), .A2(result[11]), .A3(n4980), .A4(
        result[14]), .ZN(n4074) );
  ND4D1BWP U9000 ( .A1(n3744), .A2(n3743), .A3(n3742), .A4(n3741), .ZN(
        result[14]) );
  OAI211D1BWP U9001 ( .A1(n5791), .A2(n5790), .B(n4656), .C(n5789), .ZN(
        \alu/N665 ) );
  AOI222D1BWP U9002 ( .A1(n5788), .A2(n5791), .B1(n5788), .B2(n5787), .C1(
        n5791), .C2(n5786), .ZN(n5789) );
  IND2D1BWP U9003 ( .A1(n5782), .B1(n4659), .ZN(n5783) );
  AOI21D1BWP U9004 ( .A1(n4836), .A2(n4835), .B(n4834), .ZN(\alu/N1018 ) );
  AOI32D1BWP U9005 ( .A1(n5691), .A2(n5804), .A3(n5690), .B1(n5689), .B2(n5804), .ZN(\alu/N1003 ) );
  AOI22D1BWP U9006 ( .A1(n4672), .A2(\alu/N683 ), .B1(n4671), .B2(op2[6]), 
        .ZN(n3744) );
  NR2XD0BWP U9007 ( .A1(\intadd_34/A[1] ), .A2(\intadd_34/A[2] ), .ZN(n4980)
         );
  NR2XD0BWP U9008 ( .A1(n5781), .A2(n5780), .ZN(n5787) );
  NR2XD0BWP U9009 ( .A1(n5769), .A2(n5768), .ZN(n5775) );
  NR2XD0BWP U9010 ( .A1(n5765), .A2(n5767), .ZN(n5771) );
  NR2XD0BWP U9011 ( .A1(n5774), .A2(n5773), .ZN(n5765) );
  AOI21D1BWP U9012 ( .A1(n5768), .A2(n5782), .B(n5778), .ZN(n5767) );
  NR2XD0BWP U9013 ( .A1(n5782), .A2(n5768), .ZN(n5778) );
  AOI22D1BWP U9014 ( .A1(op2[2]), .A2(n4671), .B1(\alu/N1014 ), .B2(n4690), 
        .ZN(n6066) );
  AOI22D1BWP U9015 ( .A1(n4689), .A2(\alu/N661 ), .B1(n4672), .B2(op1[10]), 
        .ZN(n6065) );
  OAI211D1BWP U9016 ( .A1(n5764), .A2(n5790), .B(n4656), .C(n5763), .ZN(
        \alu/N661 ) );
  OAI21D1BWP U9017 ( .A1(n5788), .A2(n5762), .B(n5766), .ZN(n5763) );
  AOI21D1BWP U9018 ( .A1(n5788), .A2(n5762), .B(n5761), .ZN(n5766) );
  AOI21D1BWP U9019 ( .A1(n5762), .A2(n5760), .B(n5773), .ZN(n5764) );
  NR2XD0BWP U9020 ( .A1(n5760), .A2(n5762), .ZN(n5773) );
  OAI21D1BWP U9021 ( .A1(n4465), .A2(n4464), .B(n5782), .ZN(n5769) );
  AOI22D1BWP U9022 ( .A1(n4692), .A2(\alu/N832 ), .B1(n4691), .B2(\alu/N832 ), 
        .ZN(n6064) );
  OAI31D1BWP U9023 ( .A1(n5683), .A2(n5689), .A3(n5682), .B(n5681), .ZN(n5804)
         );
  OAI21D1BWP U9024 ( .A1(n5683), .A2(n5682), .B(n5689), .ZN(n5681) );
  AOI222D1BWP U9025 ( .A1(n5680), .A2(n5679), .B1(n5680), .B2(n5678), .C1(
        n5679), .C2(n5677), .ZN(n5682) );
  IND2D1BWP U9026 ( .A1(n5676), .B1(n5675), .ZN(n5677) );
  NR2XD0BWP U9027 ( .A1(n5691), .A2(n5690), .ZN(n5689) );
  NR2XD0BWP U9028 ( .A1(n5687), .A2(n5688), .ZN(n5690) );
  OAI211D1BWP U9029 ( .A1(\intadd_36/SUM[2] ), .A2(n5672), .B(n5671), .C(n5670), .ZN(n5688) );
  OAI211D1BWP U9030 ( .A1(n5669), .A2(n5668), .B(n5667), .C(n5676), .ZN(n5670)
         );
  AOI22D1BWP U9031 ( .A1(n5666), .A2(n5669), .B1(n5665), .B2(n5664), .ZN(n5671) );
  AOI211XD0BWP U9032 ( .A1(n5661), .A2(n5665), .B(n5660), .C(n5659), .ZN(n5685) );
  OAI22D1BWP U9033 ( .A1(n5658), .A2(n5680), .B1(n5657), .B2(n5678), .ZN(n5659) );
  XNR2D1BWP U9034 ( .A1(n5657), .A2(n5656), .ZN(n5658) );
  NR2XD0BWP U9035 ( .A1(n5672), .A2(\intadd_36/SUM[1] ), .ZN(n5660) );
  NR2XD0BWP U9036 ( .A1(n5684), .A2(n5803), .ZN(n5686) );
  AO221D1BWP U9037 ( .A1(n5678), .A2(n3677), .B1(n5666), .B2(n5622), .C(n5634), 
        .Z(n5803) );
  OAI211D1BWP U9038 ( .A1(\intadd_36/SUM[0] ), .A2(n5672), .B(n5627), .C(n5626), .ZN(n5684) );
  AOI32D1BWP U9039 ( .A1(n5622), .A2(n5625), .A3(n5667), .B1(n5648), .B2(n5624), .ZN(n5627) );
  OAI21D1BWP U9040 ( .A1(n5622), .A2(n5680), .B(n5678), .ZN(n5624) );
  ND3D1BWP U9041 ( .A1(\alu/N683 ), .A2(n5795), .A3(n4658), .ZN(n5672) );
  XOR2D1BWP U9042 ( .A1(n5675), .A2(n5676), .Z(n5651) );
  NR2XD0BWP U9043 ( .A1(n5657), .A2(n5656), .ZN(n5668) );
  XNR2D1BWP U9044 ( .A1(n5674), .A2(n5645), .ZN(n5675) );
  IND2D1BWP U9045 ( .A1(n5644), .B1(n5643), .ZN(n5674) );
  AO22D1BWP U9046 ( .A1(op1[12]), .A2(n5642), .B1(n5655), .B2(n5646), .Z(n5650) );
  AOI211XD0BWP U9047 ( .A1(n4678), .A2(n5648), .B(n5641), .C(n5640), .ZN(n5642) );
  OAI22D1BWP U9048 ( .A1(n4676), .A2(n3652), .B1(n3678), .B2(op2[10]), .ZN(
        n5625) );
  OAI31D1BWP U9049 ( .A1(\alu/N684 ), .A2(n5643), .A3(\intadd_36/n1 ), .B(
        n5639), .ZN(n5653) );
  AOI21D1BWP U9050 ( .A1(n5645), .A2(n5638), .B(n5636), .ZN(n5637) );
  OAI31D1BWP U9051 ( .A1(n5638), .A2(n5636), .A3(n5673), .B(n5635), .ZN(n5683)
         );
  AOI31D1BWP U9052 ( .A1(n5643), .A2(\intadd_36/n1 ), .A3(n4658), .B(n5634), 
        .ZN(n5635) );
  IND2D1BWP U9053 ( .A1(n5640), .B1(n5630), .ZN(\intadd_36/CI ) );
  OAI21D1BWP U9054 ( .A1(op1[12]), .A2(n5640), .B(n5633), .ZN(\intadd_36/B[1] ) );
  AOI21D1BWP U9055 ( .A1(n3653), .A2(n5633), .B(n5632), .ZN(n5649) );
  OA21D1BWP U9056 ( .A1(\alu/N683 ), .A2(n5632), .B(n5704), .Z(n5643) );
  IND2D1BWP U9057 ( .A1(n5631), .B1(n5630), .ZN(n5654) );
  AOI31D1BWP U9058 ( .A1(op1[11]), .A2(n4693), .A3(n5629), .B(n5641), .ZN(
        n5631) );
  OAI21D1BWP U9059 ( .A1(op2[12]), .A2(n5641), .B(n5628), .ZN(n5647) );
  AOI21D1BWP U9060 ( .A1(n3561), .A2(n5628), .B(n4657), .ZN(n5663) );
  AOI211XD0BWP U9061 ( .A1(n4986), .A2(n4056), .B(n4055), .C(n4054), .ZN(n4642) );
  ND4D1BWP U9062 ( .A1(n4987), .A2(n6004), .A3(n6011), .A4(n6037), .ZN(n4988)
         );
  ND3D1BWP U9063 ( .A1(n6067), .A2(n6068), .A3(n6069), .ZN(result[15]) );
  AOI22D1BWP U9064 ( .A1(op2[7]), .A2(n4671), .B1(\alu/N1019 ), .B2(n4690), 
        .ZN(n6069) );
  NR2XD0BWP U9065 ( .A1(n5623), .A2(n4834), .ZN(n4986) );
  NR2XD0BWP U9066 ( .A1(n4835), .A2(n4836), .ZN(n4834) );
  MAOI222D1BWP U9067 ( .A(op1[13]), .B(op2[13]), .C(n4837), .ZN(n4836) );
  MAOI222D1BWP U9068 ( .A(n4842), .B(n4676), .C(n4677), .ZN(n4841) );
  AOI22D1BWP U9069 ( .A1(n4689), .A2(\alu/N634 ), .B1(n4672), .B2(op1[15]), 
        .ZN(n6068) );
  OAI21D1BWP U9070 ( .A1(n4692), .A2(n4691), .B(\alu/N808 ), .ZN(n6067) );
  NR2XD0BWP U9071 ( .A1(n5793), .A2(n5792), .ZN(\alu/N808 ) );
  OAI21D1BWP U9072 ( .A1(n4654), .A2(n4653), .B(n4083), .ZN(n4843) );
  OAI21D1BWP U9073 ( .A1(op1[8]), .A2(op2[8]), .B(n4846), .ZN(n4083) );
  OAI211D1BWP U9074 ( .A1(n3917), .A2(n4054), .B(n3916), .C(n3915), .ZN(
        result[8]) );
  AO22D1BWP U9075 ( .A1(n5802), .A2(\intadd_33/SUM[8] ), .B1(n5801), .B2(
        \intadd_33/SUM[7] ), .Z(\alu/N990 ) );
  AOI21D1BWP U9076 ( .A1(n4689), .A2(\alu/N659 ), .B(n3914), .ZN(n3916) );
  OAI22D1BWP U9077 ( .A1(n3913), .A2(n4653), .B1(n3912), .B2(n4680), .ZN(n3914) );
  NR2XD0BWP U9078 ( .A1(n5759), .A2(n5757), .ZN(\alu/N659 ) );
  XNR3D1BWP U9079 ( .A1(n4846), .A2(op1[8]), .A3(op2[8]), .ZN(n3917) );
  OAI21D1BWP U9080 ( .A1(n4833), .A2(n5605), .B(n4847), .ZN(n4846) );
  OAI211D1BWP U9081 ( .A1(n5755), .A2(n3901), .B(n3900), .C(n3899), .ZN(n3902)
         );
  AO22D1BWP U9082 ( .A1(n5802), .A2(\intadd_33/SUM[7] ), .B1(n5801), .B2(
        \intadd_33/SUM[6] ), .Z(\alu/N989 ) );
  AOI21D1BWP U9083 ( .A1(n4690), .A2(\alu/N1011 ), .B(n3898), .ZN(n3900) );
  OAI22D1BWP U9084 ( .A1(n3913), .A2(n4833), .B1(n3912), .B2(n5605), .ZN(n3898) );
  OA21D1BWP U9085 ( .A1(n4849), .A2(n4848), .B(n4847), .Z(\alu/N1011 ) );
  OAI21D1BWP U9086 ( .A1(n4662), .A2(n4663), .B(n4082), .ZN(n4848) );
  OAI21D1BWP U9087 ( .A1(op1[6]), .A2(op2[6]), .B(n4850), .ZN(n4082) );
  AOI211XD0BWP U9088 ( .A1(n5752), .A2(n5751), .B(n5750), .C(n5790), .ZN(n5753) );
  AOI221D1BWP U9089 ( .A1(n5774), .A2(n5746), .B1(n5745), .B2(n5744), .C(n5752), .ZN(n5750) );
  OAI32D1BWP U9090 ( .A1(n5774), .A2(n5743), .A3(n5742), .B1(n5741), .B2(n5745), .ZN(n5751) );
  AOI22D1BWP U9091 ( .A1(n5760), .A2(n5755), .B1(n5740), .B2(n5739), .ZN(n5742) );
  AOI211XD0BWP U9092 ( .A1(n5748), .A2(n5747), .B(n5738), .C(n5737), .ZN(n5743) );
  INR2D1BWP U9093 ( .A1(n5734), .B1(n5735), .ZN(n5772) );
  INR2D1BWP U9094 ( .A1(n5733), .B1(n5732), .ZN(n5735) );
  NR2XD0BWP U9095 ( .A1(n5731), .A2(n5730), .ZN(n5734) );
  MUX2ND0BWP U9096 ( .I0(n3799), .I1(n3888), .S(n4674), .ZN(n4673) );
  INR2D1BWP U9097 ( .A1(n5726), .B1(n4644), .ZN(n5747) );
  AOI21D1BWP U9098 ( .A1(n5757), .A2(n5725), .B(n5730), .ZN(n5760) );
  XOR2D1BWP U9099 ( .A1(n4624), .A2(n5724), .Z(n5730) );
  AOI32D1BWP U9100 ( .A1(n5736), .A2(n5755), .A3(n5723), .B1(n5722), .B2(n5755), .ZN(n5725) );
  AOI32D1BWP U9101 ( .A1(n5726), .A2(n5728), .A3(n4644), .B1(n5719), .B2(n5728), .ZN(n5723) );
  OAI21D1BWP U9102 ( .A1(n5718), .A2(n5717), .B(n5724), .ZN(n5757) );
  NR2XD0BWP U9103 ( .A1(n4445), .A2(n5720), .ZN(n5718) );
  XOR2D1BWP U9104 ( .A1(n5710), .A2(n5709), .Z(n5727) );
  XOR2D1BWP U9105 ( .A1(n5714), .A2(n5715), .Z(n5736) );
  OAI211D1BWP U9106 ( .A1(n3853), .A2(n4054), .B(n3852), .C(n3851), .ZN(
        result[6]) );
  AO22D1BWP U9107 ( .A1(n5802), .A2(\intadd_33/SUM[6] ), .B1(n5801), .B2(
        \intadd_33/SUM[5] ), .Z(\alu/N988 ) );
  AOI21D1BWP U9108 ( .A1(n4689), .A2(\alu/N657 ), .B(n3850), .ZN(n3852) );
  OAI22D1BWP U9109 ( .A1(n3913), .A2(n4663), .B1(n3912), .B2(n4662), .ZN(n3850) );
  NR2XD0BWP U9110 ( .A1(n5754), .A2(n5740), .ZN(\alu/N657 ) );
  XOR2D1BWP U9111 ( .A1(n5721), .A2(n5720), .Z(n5740) );
  XNR3D1BWP U9112 ( .A1(op1[6]), .A2(op2[6]), .A3(n4850), .ZN(n3853) );
  OAI21D1BWP U9113 ( .A1(n4666), .A2(n4667), .B(n4081), .ZN(n4851) );
  OAI21D1BWP U9114 ( .A1(op1[4]), .A2(op2[4]), .B(n4854), .ZN(n4081) );
  OAI211D1BWP U9115 ( .A1(n3814), .A2(n4054), .B(n3813), .C(n3812), .ZN(
        result[2]) );
  AO22D1BWP U9116 ( .A1(n5802), .A2(\intadd_33/SUM[2] ), .B1(n5801), .B2(
        \intadd_33/SUM[1] ), .Z(\alu/N984 ) );
  AOI21D1BWP U9117 ( .A1(n4689), .A2(\alu/N653 ), .B(n3811), .ZN(n3813) );
  OAI22D1BWP U9118 ( .A1(n3913), .A2(n4670), .B1(n3912), .B2(n4669), .ZN(n3811) );
  NR2XD0BWP U9119 ( .A1(n5754), .A2(n5726), .ZN(\alu/N653 ) );
  XNR2D1BWP U9120 ( .A1(n5707), .A2(n5708), .ZN(n5726) );
  XNR3D1BWP U9121 ( .A1(n4857), .A2(op2[2]), .A3(op1[2]), .ZN(n3814) );
  OAI211D1BWP U9122 ( .A1(n3837), .A2(n4054), .B(n3836), .C(n3835), .ZN(
        result[4]) );
  AO22D1BWP U9123 ( .A1(n5802), .A2(\intadd_33/SUM[4] ), .B1(n5801), .B2(
        \intadd_33/SUM[3] ), .Z(\alu/N986 ) );
  AOI21D1BWP U9124 ( .A1(n4689), .A2(\alu/N655 ), .B(n3834), .ZN(n3836) );
  OAI22D1BWP U9125 ( .A1(n3913), .A2(n4667), .B1(n3912), .B2(n4666), .ZN(n3834) );
  NR2XD0BWP U9126 ( .A1(n5754), .A2(n5728), .ZN(\alu/N655 ) );
  NR2XD0BWP U9127 ( .A1(n5712), .A2(n5711), .ZN(n5716) );
  NR2XD0BWP U9128 ( .A1(n5711), .A2(n5706), .ZN(n5708) );
  XNR3D1BWP U9129 ( .A1(op1[4]), .A2(op2[4]), .A3(n4854), .ZN(n3837) );
  OAI21D1BWP U9130 ( .A1(n4669), .A2(n4670), .B(n4080), .ZN(n4855) );
  OAI21D1BWP U9131 ( .A1(op2[2]), .A2(op1[2]), .B(n4857), .ZN(n4080) );
  NR2XD0BWP U9132 ( .A1(n4858), .A2(n4859), .ZN(n4857) );
  OAI211D1BWP U9133 ( .A1(n5729), .A2(n3901), .B(n3804), .C(n3803), .ZN(
        result[1]) );
  OAI21D1BWP U9134 ( .A1(n4672), .A2(n3802), .B(op2[1]), .ZN(n3803) );
  AOI21D1BWP U9135 ( .A1(n4860), .A2(n4701), .B(n4054), .ZN(n3802) );
  AOI21D1BWP U9136 ( .A1(\alu/N983 ), .A2(n3925), .B(n3801), .ZN(n3804) );
  OAI22D1BWP U9137 ( .A1(n4861), .A2(n4054), .B1(n3912), .B2(n6070), .ZN(n3801) );
  NR2XD0BWP U9138 ( .A1(op1[1]), .A2(n4862), .ZN(n4858) );
  NR2XD0BWP U9139 ( .A1(n4679), .A2(n4680), .ZN(n4862) );
  AO22D1BWP U9140 ( .A1(n5802), .A2(\intadd_33/SUM[1] ), .B1(
        \intadd_33/SUM[0] ), .B2(n5801), .Z(\alu/N983 ) );
  NR2XD0BWP U9141 ( .A1(n5794), .A2(n5792), .ZN(n5802) );
  AOI22D1BWP U9142 ( .A1(n5621), .A2(n5620), .B1(n5619), .B2(n5618), .ZN(n5795) );
  ND4D1BWP U9143 ( .A1(n4670), .A2(n4680), .A3(n5616), .A4(n5615), .ZN(n5617)
         );
  XOR2D1BWP U9144 ( .A1(\intadd_33/n1 ), .A2(n5611), .Z(n5794) );
  OAI22D1BWP U9145 ( .A1(n5796), .A2(n5797), .B1(n5798), .B2(n5799), .ZN(
        \intadd_33/CI ) );
  MAOI222D1BWP U9146 ( .A(n5602), .B(n5601), .C(n5600), .ZN(n5603) );
  MAOI222D1BWP U9147 ( .A(\mult_x_153/n101 ), .B(\mult_x_153/n97 ), .C(n5599), 
        .ZN(n5602) );
  MAOI222D1BWP U9148 ( .A(n5598), .B(n5597), .C(n5596), .ZN(n5599) );
  MAOI222D1BWP U9149 ( .A(n5595), .B(n5594), .C(n5593), .ZN(n5597) );
  MAOI222D1BWP U9150 ( .A(n5584), .B(n5583), .C(n5582), .ZN(n5595) );
  XNR2D1BWP U9151 ( .A1(n5578), .A2(n5577), .ZN(n5579) );
  AOI211XD0BWP U9152 ( .A1(n5576), .A2(op2[0]), .B(n5575), .C(n5574), .ZN(
        n5580) );
  AOI22D1BWP U9153 ( .A1(op2[2]), .A2(n5573), .B1(op1[1]), .B2(n4670), .ZN(
        n5574) );
  AOI22D1BWP U9154 ( .A1(op1[1]), .A2(n5616), .B1(op1[0]), .B2(op2[0]), .ZN(
        n5575) );
  AOI21D1BWP U9155 ( .A1(op2[0]), .A2(n5572), .B(\mult_x_153/n162 ), .ZN(n5581) );
  OAI21D1BWP U9156 ( .A1(n6070), .A2(n4669), .B(op1[3]), .ZN(\mult_x_153/n162 ) );
  IND2D1BWP U9157 ( .A1(n5578), .B1(n5577), .ZN(n5583) );
  OAI31D1BWP U9158 ( .A1(op1[0]), .A2(op2[2]), .A3(n6070), .B(n5571), .ZN(
        n5577) );
  AOI22D1BWP U9159 ( .A1(op2[3]), .A2(n5570), .B1(\mult_x_153/n176 ), .B2(
        n5569), .ZN(n5571) );
  OAI32D1BWP U9160 ( .A1(n4669), .A2(n4680), .A3(op1[3]), .B1(n5566), .B2(
        op2[0]), .ZN(n5568) );
  AOI21D1BWP U9161 ( .A1(op2[4]), .A2(n5570), .B(n5565), .ZN(n5585) );
  OAI22D1BWP U9162 ( .A1(op2[3]), .A2(n5564), .B1(op2[4]), .B2(n5573), .ZN(
        n5565) );
  AOI22D1BWP U9163 ( .A1(op1[3]), .A2(n5616), .B1(op2[1]), .B2(n5561), .ZN(
        n5567) );
  AO21D1BWP U9164 ( .A1(n5560), .A2(n5559), .B(\mult_x_153/n105 ), .Z(n5589)
         );
  AOI21D1BWP U9165 ( .A1(op2[5]), .A2(n5570), .B(n5558), .ZN(n5590) );
  OAI22D1BWP U9166 ( .A1(op2[5]), .A2(n5573), .B1(op2[4]), .B2(n5564), .ZN(
        n5558) );
  AOI22D1BWP U9167 ( .A1(n5563), .A2(n5557), .B1(n5556), .B2(n5572), .ZN(n5591) );
  OAI22D1BWP U9168 ( .A1(n5561), .A2(n5569), .B1(op2[3]), .B2(op1[3]), .ZN(
        n4856) );
  AOI22D1BWP U9169 ( .A1(op1[3]), .A2(op2[2]), .B1(n4670), .B2(n5561), .ZN(
        n5563) );
  OAI32D1BWP U9170 ( .A1(op1[9]), .A2(n5555), .A3(n4653), .B1(n5554), .B2(
        n3680), .ZN(n5607) );
  OAI21D1BWP U9171 ( .A1(n5606), .A2(n5608), .B(n5609), .ZN(\intadd_33/A[9] )
         );
  AOI22D1BWP U9172 ( .A1(op1[9]), .A2(op2[8]), .B1(op2[9]), .B2(n3680), .ZN(
        n5608) );
  OA31D1BWP U9173 ( .A1(n4653), .A2(n5605), .A3(n4648), .B(n5610), .Z(n5606)
         );
  AOI21D1BWP U9174 ( .A1(n4648), .A2(n5604), .B(n3680), .ZN(n5610) );
  NR2XD0BWP U9175 ( .A1(n5788), .A2(n5761), .ZN(n5786) );
  IND3D1BWP U9176 ( .A1(n4457), .B1(n4456), .B2(n4455), .ZN(n5756) );
  NR2XD0BWP U9177 ( .A1(n5724), .A2(n4624), .ZN(n5788) );
  NR2XD0BWP U9178 ( .A1(n3561), .A2(n5628), .ZN(n4657) );
  NR2XD0BWP U9179 ( .A1(n4693), .A2(n4676), .ZN(n5641) );
  OAI21D1BWP U9180 ( .A1(n3896), .A2(n4411), .B(n3895), .ZN(n4464) );
  MUX2ND0BWP U9181 ( .I0(n3894), .I1(\alu/N339 ), .S(n4675), .ZN(n3895) );
  AOI21D1BWP U9182 ( .A1(n4449), .A2(n3893), .B(\intadd_35/CI ), .ZN(n3896) );
  NR4D0BWP U9183 ( .A1(n5700), .A2(n5701), .A3(n3892), .A4(n3891), .ZN(n4463)
         );
  XOR2D1BWP U9184 ( .A1(n3890), .A2(n3889), .Z(n3891) );
  XOR2D1BWP U9185 ( .A1(n3799), .A2(n3800), .Z(n3888) );
  OAI221D1BWP U9186 ( .A1(n5710), .A2(n5697), .B1(n5706), .B2(n5707), .C(n5696), .ZN(n5701) );
  AOI22D1BWP U9187 ( .A1(n5697), .A2(n5707), .B1(n5706), .B2(n5710), .ZN(n5696) );
  NR4D0BWP U9188 ( .A1(n5721), .A2(n4446), .A3(n5715), .A4(n5717), .ZN(n5698)
         );
  ND4D1BWP U9189 ( .A1(n4645), .A2(n5713), .A3(n5707), .A4(n5710), .ZN(n5712)
         );
  AO21D1BWP U9190 ( .A1(n4441), .A2(n4427), .B(n4426), .Z(n5710) );
  OAI31D1BWP U9191 ( .A1(\intadd_35/B[0] ), .A2(n4425), .A3(n4444), .B(n4424), 
        .ZN(n4426) );
  AOI22D1BWP U9192 ( .A1(\alu/N339 ), .A2(\alu/N332 ), .B1(\alu/N331 ), .B2(
        n4451), .ZN(n4424) );
  AO222D1BWP U9193 ( .A1(n4451), .A2(\alu/N330 ), .B1(n4423), .B2(n4422), .C1(
        \alu/N331 ), .C2(\alu/N339 ), .Z(n5707) );
  OAI21D1BWP U9194 ( .A1(n4421), .A2(n4444), .B(n4420), .ZN(n4422) );
  ND3D1BWP U9195 ( .A1(n4457), .A2(n4455), .A3(n4419), .ZN(n4420) );
  OAI211D1BWP U9196 ( .A1(n4444), .A2(n4437), .B(n4418), .C(n4417), .ZN(n5713)
         );
  AOI22D1BWP U9197 ( .A1(\alu/N339 ), .A2(\alu/N333 ), .B1(\alu/N332 ), .B2(
        n4451), .ZN(n4418) );
  OAI211D1BWP U9198 ( .A1(n4448), .A2(n4437), .B(n4436), .C(n4435), .ZN(n5717)
         );
  MUX2ND0BWP U9199 ( .I0(n4416), .I1(n4415), .S(\intadd_35/B[0] ), .ZN(n4434)
         );
  AOI21D1BWP U9200 ( .A1(n4433), .A2(n4432), .B(n4431), .ZN(n4436) );
  AOI21D1BWP U9201 ( .A1(\alu/N335 ), .A2(n4428), .B(\alu/N339 ), .ZN(n4430)
         );
  OAI211D1BWP U9202 ( .A1(n4444), .A2(n4447), .B(n4443), .C(n4442), .ZN(n5715)
         );
  MUX2ND0BWP U9203 ( .I0(n4440), .I1(n4439), .S(\intadd_35/B[0] ), .ZN(n4454)
         );
  AOI22D1BWP U9204 ( .A1(\alu/N339 ), .A2(\alu/N334 ), .B1(\alu/N333 ), .B2(
        n4451), .ZN(n4443) );
  MUX2ND0BWP U9205 ( .I0(\alu/N332 ), .I1(\alu/N333 ), .S(n4449), .ZN(n4440)
         );
  MUX2ND0BWP U9206 ( .I0(n4439), .I1(n3882), .S(\intadd_35/B[0] ), .ZN(n4427)
         );
  MUX2ND0BWP U9207 ( .I0(\alu/N330 ), .I1(\alu/N331 ), .S(n4449), .ZN(n4439)
         );
  OAI211D1BWP U9208 ( .A1(n4416), .A2(n4452), .B(n3881), .C(n3880), .ZN(n5721)
         );
  NR2XD0BWP U9209 ( .A1(n4419), .A2(n4410), .ZN(n4453) );
  MUX2ND0BWP U9210 ( .I0(n4415), .I1(n3879), .S(\intadd_35/B[0] ), .ZN(n4457)
         );
  MUX2ND0BWP U9211 ( .I0(\alu/N329 ), .I1(\alu/N330 ), .S(n4449), .ZN(n4415)
         );
  AOI31D1BWP U9212 ( .A1(n4441), .A2(n3878), .A3(n4432), .B(n3877), .ZN(n3881)
         );
  OAI21D1BWP U9213 ( .A1(n4448), .A2(n4421), .B(n3876), .ZN(n3877) );
  AOI22D1BWP U9214 ( .A1(\alu/N339 ), .A2(\alu/N335 ), .B1(\alu/N334 ), .B2(
        n4451), .ZN(n3876) );
  ND3D1BWP U9215 ( .A1(\alu/N326 ), .A2(n3875), .A3(n3874), .ZN(n4421) );
  MUX2ND0BWP U9216 ( .I0(n3873), .I1(n3872), .S(n4449), .ZN(n4432) );
  MUX2ND0BWP U9217 ( .I0(\alu/N331 ), .I1(\alu/N332 ), .S(n4449), .ZN(n4416)
         );
  NR3D0BWP U9218 ( .A1(n5780), .A2(n5770), .A3(n5768), .ZN(n4659) );
  NR2XD0BWP U9219 ( .A1(n3887), .A2(n3886), .ZN(n5768) );
  AOI211XD0BWP U9220 ( .A1(n4675), .A2(\intadd_35/A[0] ), .B(n5703), .C(n3885), 
        .ZN(n3886) );
  OAI22D1BWP U9221 ( .A1(\intadd_35/A[0] ), .A2(n3884), .B1(\intadd_35/SUM[0] ), .B2(n4411), .ZN(n3887) );
  OAI22D1BWP U9222 ( .A1(n5702), .A2(n3868), .B1(\intadd_35/SUM[2] ), .B2(
        n4411), .ZN(n5779) );
  OA21D1BWP U9223 ( .A1(n4455), .A2(\intadd_35/A[2] ), .B(n3869), .Z(n3868) );
  AOI21D1BWP U9224 ( .A1(n5702), .A2(n5695), .B(n5694), .ZN(n5784) );
  OAI22D1BWP U9225 ( .A1(n5702), .A2(n4413), .B1(n4412), .B2(n4411), .ZN(n5694) );
  XNR2D1BWP U9226 ( .A1(\intadd_35/n1 ), .A2(n5693), .ZN(n4412) );
  NR2XD0BWP U9227 ( .A1(n3893), .A2(n4449), .ZN(\intadd_35/CI ) );
  NR2XD0BWP U9228 ( .A1(n4423), .A2(n3864), .ZN(\intadd_35/B[2] ) );
  NR2XD0BWP U9229 ( .A1(n3869), .A2(\intadd_35/A[2] ), .ZN(n5702) );
  NR2XD0BWP U9230 ( .A1(n4675), .A2(\intadd_35/A[0] ), .ZN(n5703) );
  NR2XD0BWP U9231 ( .A1(n5633), .A2(n3653), .ZN(n5632) );
  NR2XD0BWP U9232 ( .A1(n4678), .A2(n4677), .ZN(n5640) );
  NR2XD0BWP U9233 ( .A1(n3889), .A2(n3890), .ZN(n4645) );
  MUX2ND0BWP U9234 ( .I0(op2[11]), .I1(op1[11]), .S(n4650), .ZN(
        \intadd_35/A[0] ) );
  MUX2ND0BWP U9235 ( .I0(op2[13]), .I1(op1[13]), .S(n4650), .ZN(
        \intadd_35/A[2] ) );
  MUX2ND0BWP U9236 ( .I0(op2[12]), .I1(op1[12]), .S(n4650), .ZN(
        \intadd_35/A[1] ) );
  MUX2ND0BWP U9237 ( .I0(op2[10]), .I1(op1[10]), .S(n4650), .ZN(n4675) );
  AOI31D1BWP U9238 ( .A1(n3799), .A2(n3779), .A3(n3778), .B(n4461), .ZN(n3897)
         );
  NR4D0BWP U9239 ( .A1(\alu/N321 ), .A2(\alu/N324 ), .A3(\alu/N323 ), .A4(
        \alu/N325 ), .ZN(n3774) );
  NR4D0BWP U9240 ( .A1(\alu/N317 ), .A2(\alu/N320 ), .A3(\alu/N319 ), .A4(
        \alu/N322 ), .ZN(n3775) );
  NR4D0BWP U9241 ( .A1(\alu/N314 ), .A2(\alu/N316 ), .A3(\alu/N315 ), .A4(
        \alu/N318 ), .ZN(n3776) );
  AOI222D1BWP U9242 ( .A1(\alu/N329 ), .A2(\alu/N339 ), .B1(\alu/N328 ), .B2(
        n3894), .C1(n4414), .C2(n4441), .ZN(n3799) );
  MUX2ND0BWP U9243 ( .I0(n3879), .I1(n3765), .S(\intadd_35/B[0] ), .ZN(n4414)
         );
  MUX2ND0BWP U9244 ( .I0(\alu/N327 ), .I1(\alu/N328 ), .S(n4449), .ZN(n3879)
         );
  NR2XD0BWP U9245 ( .A1(n4462), .A2(n4461), .ZN(n3800) );
  AOI222D1BWP U9246 ( .A1(n3798), .A2(n4450), .B1(\alu/N339 ), .B2(\alu/N328 ), 
        .C1(n4451), .C2(\alu/N327 ), .ZN(n4461) );
  NR2XD0BWP U9247 ( .A1(n4429), .A2(n4410), .ZN(n4450) );
  AOI22D1BWP U9248 ( .A1(\alu/N326 ), .A2(n4451), .B1(\alu/N339 ), .B2(
        \alu/N327 ), .ZN(n3779) );
  NR4D0BWP U9249 ( .A1(n3777), .A2(n3769), .A3(n3768), .A4(n3767), .ZN(n4458)
         );
  ND4D1BWP U9250 ( .A1(\alu/N321 ), .A2(\alu/N324 ), .A3(\alu/N323 ), .A4(
        \alu/N325 ), .ZN(n3767) );
  XOR2D1BWP U9251 ( .A1(\DP_OP_493J11_130_7648/n15 ), .A2(
        \DP_OP_493J11_130_7648/n44 ), .Z(\alu/N325 ) );
  XOR2D1BWP U9252 ( .A1(\DP_OP_493J11_130_7648/n17 ), .A2(
        \DP_OP_493J11_130_7648/n46 ), .Z(\alu/N323 ) );
  XOR2D1BWP U9253 ( .A1(\DP_OP_493J11_130_7648/n16 ), .A2(
        \DP_OP_493J11_130_7648/n45 ), .Z(\alu/N324 ) );
  XOR2D1BWP U9254 ( .A1(\DP_OP_493J11_130_7648/n19 ), .A2(
        \DP_OP_493J11_130_7648/n48 ), .Z(\alu/N321 ) );
  ND4D1BWP U9255 ( .A1(\alu/N317 ), .A2(\alu/N320 ), .A3(\alu/N319 ), .A4(
        \alu/N322 ), .ZN(n3768) );
  XOR2D1BWP U9256 ( .A1(\DP_OP_493J11_130_7648/n18 ), .A2(
        \DP_OP_493J11_130_7648/n47 ), .Z(\alu/N322 ) );
  XOR2D1BWP U9257 ( .A1(\DP_OP_493J11_130_7648/n21 ), .A2(
        \DP_OP_493J11_130_7648/n50 ), .Z(\alu/N319 ) );
  XOR2D1BWP U9258 ( .A1(\DP_OP_493J11_130_7648/n20 ), .A2(
        \DP_OP_493J11_130_7648/n49 ), .Z(\alu/N320 ) );
  XOR2D1BWP U9259 ( .A1(\DP_OP_493J11_130_7648/n23 ), .A2(
        \DP_OP_493J11_130_7648/n52 ), .Z(\alu/N317 ) );
  ND4D1BWP U9260 ( .A1(\alu/N314 ), .A2(\alu/N316 ), .A3(\alu/N315 ), .A4(
        \alu/N318 ), .ZN(n3769) );
  XOR2D1BWP U9261 ( .A1(\DP_OP_493J11_130_7648/n22 ), .A2(
        \DP_OP_493J11_130_7648/n51 ), .Z(\alu/N318 ) );
  XOR2D1BWP U9262 ( .A1(\DP_OP_493J11_130_7648/n25 ), .A2(
        \DP_OP_493J11_130_7648/n54 ), .Z(\alu/N315 ) );
  XOR2D1BWP U9263 ( .A1(\DP_OP_493J11_130_7648/n24 ), .A2(
        \DP_OP_493J11_130_7648/n53 ), .Z(\alu/N316 ) );
  XOR2D1BWP U9264 ( .A1(\DP_OP_493J11_130_7648/n26 ), .A2(
        \DP_OP_493J11_130_7648/n55 ), .Z(\alu/N314 ) );
  MUX2ND0BWP U9265 ( .I0(\alu/N313 ), .I1(\alu/N326 ), .S(\alu/N339 ), .ZN(
        n3777) );
  XOR2D1BWP U9266 ( .A1(\DP_OP_493J11_130_7648/n56 ), .A2(n4612), .Z(
        \alu/N313 ) );
  AOI222D1BWP U9267 ( .A1(n4451), .A2(\alu/N329 ), .B1(\alu/N339 ), .B2(
        \alu/N330 ), .C1(n4441), .C2(n4438), .ZN(n3890) );
  MUX2ND0BWP U9268 ( .I0(n3882), .I1(n4425), .S(\intadd_35/B[0] ), .ZN(n4438)
         );
  AOI21D1BWP U9269 ( .A1(n3766), .A2(n3874), .B(\alu/N337 ), .ZN(
        \intadd_35/B[0] ) );
  IOA21D1BWP U9270 ( .A1(\alu/N328 ), .A2(n3773), .B(n3770), .ZN(n3764) );
  MUX2D1BWP U9271 ( .I0(\alu/N326 ), .I1(\alu/N327 ), .S(n4449), .Z(n3798) );
  XOR2D1BWP U9272 ( .A1(\DP_OP_493J11_130_7648/n13 ), .A2(
        \DP_OP_493J11_130_7648/n42 ), .Z(\alu/N327 ) );
  MUX2ND0BWP U9273 ( .I0(\alu/N328 ), .I1(\alu/N329 ), .S(n4449), .ZN(n3882)
         );
  NR2XD0BWP U9274 ( .A1(n3763), .A2(\alu/N337 ), .ZN(n4449) );
  NR2XD0BWP U9275 ( .A1(\alu/N336 ), .A2(n3762), .ZN(n3763) );
  AOI21D1BWP U9276 ( .A1(n3872), .A2(n3761), .B(\alu/N335 ), .ZN(n3762) );
  OAI21D1BWP U9277 ( .A1(\alu/N332 ), .A2(n3760), .B(n3873), .ZN(n3761) );
  AOI21D1BWP U9278 ( .A1(\alu/N329 ), .A2(n3759), .B(\alu/N331 ), .ZN(n3760)
         );
  NR2XD0BWP U9279 ( .A1(n4410), .A2(n3772), .ZN(n4441) );
  OAI21D1BWP U9280 ( .A1(\alu/N339 ), .A2(n3867), .B(n3884), .ZN(n4451) );
  NR2XD0BWP U9281 ( .A1(n4428), .A2(\alu/N339 ), .ZN(n3894) );
  NR2XD0BWP U9282 ( .A1(\alu/N330 ), .A2(\alu/N329 ), .ZN(n3773) );
  NR2XD0BWP U9283 ( .A1(n3865), .A2(n3866), .ZN(n4456) );
  NR2XD0BWP U9284 ( .A1(\alu/N336 ), .A2(\alu/N335 ), .ZN(n3766) );
  NR2XD0BWP U9285 ( .A1(\alu/N332 ), .A2(\alu/N331 ), .ZN(n3770) );
  NR2XD0BWP U9286 ( .A1(\alu/N334 ), .A2(\alu/N333 ), .ZN(n3771) );
  NR2XD0BWP U9287 ( .A1(n3658), .A2(n3659), .ZN(\DP_OP_493J11_130_7648/n12 )
         );
  MUX2ND0BWP U9288 ( .I0(n3981), .I1(n3980), .S(n4650), .ZN(n4589) );
  AOI222D1BWP U9289 ( .A1(n3619), .A2(n4002), .B1(n3989), .B2(n4035), .C1(
        n4013), .C2(n4023), .ZN(n3980) );
  AOI222D1BWP U9290 ( .A1(n3618), .A2(n4002), .B1(n3989), .B2(n4032), .C1(
        n4011), .C2(n4023), .ZN(n3981) );
  MUX2ND0BWP U9291 ( .I0(n3985), .I1(n3984), .S(n4650), .ZN(n4588) );
  AOI222D1BWP U9292 ( .A1(n4019), .A2(n4002), .B1(n4754), .B2(n3989), .C1(
        n4018), .C2(n4003), .ZN(n3984) );
  AOI222D1BWP U9293 ( .A1(n4017), .A2(n4002), .B1(n4732), .B2(n3989), .C1(
        n4016), .C2(n4003), .ZN(n3985) );
  MUX2ND0BWP U9294 ( .I0(n3991), .I1(n3990), .S(n4650), .ZN(n4587) );
  AOI222D1BWP U9295 ( .A1(n4024), .A2(n4003), .B1(n3989), .B2(n4047), .C1(
        n4002), .C2(n4741), .ZN(n3990) );
  AOI222D1BWP U9296 ( .A1(n4022), .A2(n4003), .B1(n3989), .B2(n4045), .C1(
        n4002), .C2(n4720), .ZN(n3991) );
  MUX2ND0BWP U9297 ( .I0(n3995), .I1(n3994), .S(n4650), .ZN(n4586) );
  AOI22D1BWP U9298 ( .A1(n4002), .A2(n4748), .B1(n4003), .B2(n4028), .ZN(n3994) );
  AOI22D1BWP U9299 ( .A1(n4728), .A2(n4002), .B1(n4003), .B2(n4027), .ZN(n3995) );
  MUX2ND0BWP U9300 ( .I0(n3997), .I1(n3996), .S(n4650), .ZN(n4585) );
  MUX2ND0BWP U9301 ( .I0(n4001), .I1(n4000), .S(n4650), .ZN(n4584) );
  AOI222D1BWP U9302 ( .A1(n4002), .A2(n4754), .B1(n4003), .B2(n4756), .C1(
        n4049), .C2(n4040), .ZN(n4000) );
  AOI222D1BWP U9303 ( .A1(n4002), .A2(n4732), .B1(n4003), .B2(n4734), .C1(
        n4049), .C2(n4039), .ZN(n4001) );
  MUX2ND0BWP U9304 ( .I0(n4005), .I1(n4004), .S(n4650), .ZN(n4583) );
  AOI222D1BWP U9305 ( .A1(n4051), .A2(n4012), .B1(n4003), .B2(n4755), .C1(
        n4002), .C2(n4047), .ZN(n4004) );
  AOI222D1BWP U9306 ( .A1(n4046), .A2(n4012), .B1(n4003), .B2(n4733), .C1(
        n4002), .C2(n4045), .ZN(n4005) );
  MUX2ND0BWP U9307 ( .I0(n4010), .I1(n4009), .S(n4650), .ZN(n4582) );
  AOI222D1BWP U9308 ( .A1(n4748), .A2(n4023), .B1(n4749), .B2(n4048), .C1(
        n4008), .C2(n4012), .ZN(n4009) );
  AOI222D1BWP U9309 ( .A1(n4728), .A2(n4023), .B1(n4729), .B2(n4048), .C1(
        n4007), .C2(n4012), .ZN(n4010) );
  MUX2ND0BWP U9310 ( .I0(n4015), .I1(n4014), .S(n4650), .ZN(n4581) );
  AOI222D1BWP U9311 ( .A1(n3619), .A2(n4048), .B1(n4023), .B2(n4035), .C1(
        n4013), .C2(n4012), .ZN(n4014) );
  AOI222D1BWP U9312 ( .A1(n3618), .A2(n4048), .B1(n4023), .B2(n4032), .C1(
        n4011), .C2(n4012), .ZN(n4015) );
  NR2XD0BWP U9313 ( .A1(n4034), .A2(n4649), .ZN(n4012) );
  MUX2ND0BWP U9314 ( .I0(n4021), .I1(n4020), .S(n4650), .ZN(n4580) );
  AOI222D1BWP U9315 ( .A1(n4019), .A2(n4048), .B1(n4754), .B2(n4023), .C1(
        n4018), .C2(n4049), .ZN(n4020) );
  AOI222D1BWP U9316 ( .A1(n4017), .A2(n4048), .B1(n4732), .B2(n4023), .C1(
        n4016), .C2(n4049), .ZN(n4021) );
  MUX2ND0BWP U9317 ( .I0(n4026), .I1(n4025), .S(n4650), .ZN(n4579) );
  AOI222D1BWP U9318 ( .A1(n4024), .A2(n4049), .B1(n4047), .B2(n4023), .C1(
        n4048), .C2(n4741), .ZN(n4025) );
  AOI222D1BWP U9319 ( .A1(n4022), .A2(n4049), .B1(n4045), .B2(n4023), .C1(
        n4048), .C2(n4720), .ZN(n4026) );
  MUX2ND0BWP U9320 ( .I0(n4030), .I1(n4029), .S(n4650), .ZN(n4578) );
  AOI22D1BWP U9321 ( .A1(n4748), .A2(n4048), .B1(n4028), .B2(n4049), .ZN(n4029) );
  AOI22D1BWP U9322 ( .A1(n4728), .A2(n4048), .B1(n4027), .B2(n4049), .ZN(n4030) );
  MUX2ND0BWP U9323 ( .I0(n4037), .I1(n4036), .S(n4650), .ZN(n4577) );
  MUX2ND0BWP U9324 ( .I0(n4739), .I1(n3979), .S(n3678), .ZN(n4035) );
  MUX2ND0BWP U9325 ( .I0(n4719), .I1(n3978), .S(n3678), .ZN(n4032) );
  MUX2ND0BWP U9326 ( .I0(n4042), .I1(n4041), .S(n4650), .ZN(n4576) );
  AOI222D1BWP U9327 ( .A1(n4048), .A2(n4754), .B1(n4049), .B2(n4756), .C1(
        n4040), .C2(n4043), .ZN(n4041) );
  NR2XD0BWP U9328 ( .A1(n3678), .A2(n4744), .ZN(n4754) );
  AOI222D1BWP U9329 ( .A1(n4048), .A2(n4732), .B1(n4049), .B2(n4734), .C1(
        n4039), .C2(n4043), .ZN(n4042) );
  NR2XD0BWP U9330 ( .A1(n3678), .A2(n4724), .ZN(n4732) );
  MUX2ND0BWP U9331 ( .I0(n4053), .I1(n4052), .S(n4650), .ZN(n4575) );
  AOI222D1BWP U9332 ( .A1(n4051), .A2(n4050), .B1(n4049), .B2(n4755), .C1(
        n4048), .C2(n4047), .ZN(n4052) );
  NR2XD0BWP U9333 ( .A1(n3988), .A2(n4680), .ZN(n4047) );
  AOI222D1BWP U9334 ( .A1(n4046), .A2(n4050), .B1(n4049), .B2(n4733), .C1(
        n4048), .C2(n4045), .ZN(n4053) );
  NR2XD0BWP U9335 ( .A1(n3988), .A2(n4679), .ZN(n4045) );
  NR2XD0BWP U9336 ( .A1(n4006), .A2(n4751), .ZN(n4048) );
  NR2XD0BWP U9337 ( .A1(n3999), .A2(n4038), .ZN(n4049) );
  NR2XD0BWP U9338 ( .A1(n4044), .A2(n4649), .ZN(n4050) );
  NR2XD0BWP U9339 ( .A1(n4038), .A2(n4753), .ZN(n4043) );
  MUX2ND0BWP U9340 ( .I0(n4680), .I1(n4679), .S(n4650), .ZN(n4601) );
  MUX2ND0BWP U9341 ( .I0(n3977), .I1(n3976), .S(n4650), .ZN(n4590) );
  AOI222D1BWP U9342 ( .A1(n4002), .A2(n4749), .B1(n4748), .B2(n3989), .C1(
        n4008), .C2(n4023), .ZN(n3976) );
  AOI22D1BWP U9343 ( .A1(n3652), .A2(n4745), .B1(n4744), .B2(n3678), .ZN(n4748) );
  AOI22D1BWP U9344 ( .A1(n5622), .A2(op2[1]), .B1(op2[0]), .B2(n3677), .ZN(
        n4744) );
  AOI222D1BWP U9345 ( .A1(n4728), .A2(n3989), .B1(n4002), .B2(n4729), .C1(
        n4007), .C2(n4023), .ZN(n3977) );
  NR2XD0BWP U9346 ( .A1(n3975), .A2(n4751), .ZN(n4002) );
  AOI22D1BWP U9347 ( .A1(n3652), .A2(n4725), .B1(n4724), .B2(n3678), .ZN(n4728) );
  AOI22D1BWP U9348 ( .A1(n5622), .A2(op1[1]), .B1(op1[0]), .B2(n3677), .ZN(
        n4724) );
  MUX2ND0BWP U9349 ( .I0(n5616), .I1(n6070), .S(n4650), .ZN(n4602) );
  MUX2ND0BWP U9350 ( .I0(n3974), .I1(n3973), .S(n4650), .ZN(n4591) );
  AOI22D1BWP U9351 ( .A1(n3972), .A2(n4755), .B1(n4023), .B2(n4051), .ZN(n3973) );
  OAI22D1BWP U9352 ( .A1(n3677), .A2(op2[2]), .B1(op2[1]), .B2(n5622), .ZN(
        n4739) );
  AOI22D1BWP U9353 ( .A1(n3972), .A2(n4733), .B1(n4023), .B2(n4046), .ZN(n3974) );
  NR2XD0BWP U9354 ( .A1(n4006), .A2(n4649), .ZN(n4023) );
  OAI22D1BWP U9355 ( .A1(n3677), .A2(op1[2]), .B1(op1[1]), .B2(n5622), .ZN(
        n4719) );
  MUX2ND0BWP U9356 ( .I0(n4670), .I1(n4669), .S(n4650), .ZN(n4603) );
  MUX2ND0BWP U9357 ( .I0(n3971), .I1(n3970), .S(n4650), .ZN(n4592) );
  AOI22D1BWP U9358 ( .A1(n3972), .A2(n4756), .B1(n4003), .B2(n4040), .ZN(n3970) );
  OAI22D1BWP U9359 ( .A1(n3677), .A2(op2[3]), .B1(op2[2]), .B2(n5622), .ZN(
        n4745) );
  AOI22D1BWP U9360 ( .A1(n3972), .A2(n4734), .B1(n4003), .B2(n4039), .ZN(n3971) );
  NR2XD0BWP U9361 ( .A1(n3998), .A2(n4753), .ZN(n4003) );
  OAI22D1BWP U9362 ( .A1(n3677), .A2(op1[3]), .B1(op1[2]), .B2(n5622), .ZN(
        n4725) );
  MUX2ND0BWP U9363 ( .I0(n5569), .I1(n5561), .S(n4650), .ZN(n4604) );
  OAI22D1BWP U9364 ( .A1(n3967), .A2(n4031), .B1(n3966), .B2(n4033), .ZN(n4593) );
  MUX2ND0BWP U9365 ( .I0(n3619), .I1(n4013), .S(n4649), .ZN(n4033) );
  AOI22D1BWP U9366 ( .A1(n5622), .A2(n4667), .B1(n5569), .B2(n3677), .ZN(n4737) );
  MUX2ND0BWP U9367 ( .I0(n3618), .I1(n4011), .S(n4649), .ZN(n4031) );
  AOI22D1BWP U9368 ( .A1(n5622), .A2(n4666), .B1(n5561), .B2(n3677), .ZN(n4717) );
  MUX2ND0BWP U9369 ( .I0(n4667), .I1(n4666), .S(n4650), .ZN(n4605) );
  OAI22D1BWP U9370 ( .A1(n3992), .A2(n3967), .B1(n3993), .B2(n3966), .ZN(n4594) );
  MUX2ND0BWP U9371 ( .I0(n4749), .I1(n4008), .S(n4649), .ZN(n3993) );
  MUX2D1BWP U9372 ( .I0(n4742), .I1(n4746), .S(n3678), .Z(n4749) );
  AOI22D1BWP U9373 ( .A1(n5622), .A2(n5615), .B1(n4667), .B2(n3677), .ZN(n4746) );
  MUX2ND0BWP U9374 ( .I0(n4729), .I1(n4007), .S(n4649), .ZN(n3992) );
  MUX2D1BWP U9375 ( .I0(n4722), .I1(n4726), .S(n3678), .Z(n4729) );
  AOI22D1BWP U9376 ( .A1(n5622), .A2(n4832), .B1(n4666), .B2(n3677), .ZN(n4726) );
  MUX2ND0BWP U9377 ( .I0(n5615), .I1(n4832), .S(n4650), .ZN(n4606) );
  OAI22D1BWP U9378 ( .A1(n3987), .A2(n3966), .B1(n3986), .B2(n3967), .ZN(n4595) );
  AOI31D1BWP U9379 ( .A1(n3678), .A2(n4649), .A3(n4646), .B(n3965), .ZN(n3986)
         );
  NR2XD0BWP U9380 ( .A1(n4649), .A2(n4721), .ZN(n3965) );
  AOI22D1BWP U9381 ( .A1(n3652), .A2(n4716), .B1(n4718), .B2(n3678), .ZN(n4721) );
  AOI22D1BWP U9382 ( .A1(n5622), .A2(n4662), .B1(n4832), .B2(n3677), .ZN(n4718) );
  AOI31D1BWP U9383 ( .A1(n3678), .A2(n4649), .A3(n4647), .B(n3963), .ZN(n3987)
         );
  NR2XD0BWP U9384 ( .A1(n4649), .A2(n4740), .ZN(n3963) );
  AOI22D1BWP U9385 ( .A1(n3652), .A2(n4736), .B1(n4738), .B2(n3678), .ZN(n4740) );
  AOI22D1BWP U9386 ( .A1(n5622), .A2(n4663), .B1(n5615), .B2(n3677), .ZN(n4738) );
  MUX2ND0BWP U9387 ( .I0(n4663), .I1(n4662), .S(n4650), .ZN(n4607) );
  OAI22D1BWP U9388 ( .A1(n3983), .A2(n3966), .B1(n3982), .B2(n3967), .ZN(n4596) );
  AOI22D1BWP U9389 ( .A1(n5622), .A2(n5605), .B1(n4662), .B2(n3677), .ZN(n4722) );
  AOI22D1BWP U9390 ( .A1(n5622), .A2(n4833), .B1(n4663), .B2(n3677), .ZN(n4742) );
  MUX2ND0BWP U9391 ( .I0(n4833), .I1(n5605), .S(n4650), .ZN(n4608) );
  OAI22D1BWP U9392 ( .A1(n4747), .A2(n3958), .B1(n4727), .B2(n3957), .ZN(n4597) );
  AOI22D1BWP U9393 ( .A1(n3652), .A2(n4646), .B1(n4716), .B2(n3678), .ZN(n4727) );
  AOI22D1BWP U9394 ( .A1(n5622), .A2(n4653), .B1(n5605), .B2(n3677), .ZN(n4716) );
  AOI22D1BWP U9395 ( .A1(n3652), .A2(n4647), .B1(n4736), .B2(n3678), .ZN(n4747) );
  AOI22D1BWP U9396 ( .A1(n5622), .A2(n4654), .B1(n4833), .B2(n3677), .ZN(n4736) );
  MUX2ND0BWP U9397 ( .I0(n4654), .I1(n4653), .S(n4650), .ZN(n4609) );
  OAI22D1BWP U9398 ( .A1(n3956), .A2(n3957), .B1(n3955), .B2(n3958), .ZN(n4598) );
  MUX2ND0BWP U9399 ( .I0(n3954), .I1(n4743), .S(n3678), .ZN(n4008) );
  OAI22D1BWP U9400 ( .A1(n3677), .A2(op2[9]), .B1(op2[8]), .B2(n5622), .ZN(
        n4743) );
  MUX2ND0BWP U9401 ( .I0(n3953), .I1(n4723), .S(n3678), .ZN(n4007) );
  OAI22D1BWP U9402 ( .A1(n3677), .A2(op1[9]), .B1(op1[8]), .B2(n5622), .ZN(
        n4723) );
  MUX2ND0BWP U9403 ( .I0(n4648), .I1(n3680), .S(n4650), .ZN(n4610) );
  OAI22D1BWP U9404 ( .A1(n4735), .A2(n3958), .B1(n4715), .B2(n3957), .ZN(n4599) );
  AOI22D1BWP U9405 ( .A1(op2[10]), .A2(n3964), .B1(n3680), .B2(n3677), .ZN(
        n4646) );
  NR2XD0BWP U9406 ( .A1(n3975), .A2(n4649), .ZN(n3989) );
  AOI22D1BWP U9407 ( .A1(op1[10]), .A2(n3962), .B1(n3677), .B2(n4648), .ZN(
        n4647) );
  MUX2ND0BWP U9408 ( .I0(n3962), .I1(n3964), .S(n4650), .ZN(n4611) );
  OAI22D1BWP U9409 ( .A1(n3968), .A2(n3967), .B1(n3969), .B2(n3966), .ZN(n4600) );
  ND4D1BWP U9410 ( .A1(n3942), .A2(n4676), .A3(n4077), .A4(n4693), .ZN(
        \alu/N88 ) );
  NR2XD0BWP U9411 ( .A1(op2[13]), .A2(\alu/N684 ), .ZN(n3942) );
  OAI22D1BWP U9412 ( .A1(\alu/N683 ), .A2(n4658), .B1(n3951), .B2(n3780), .ZN(
        n5692) );
  NR2XD0BWP U9413 ( .A1(n4640), .A2(\alu/N684 ), .ZN(n3780) );
  NR2XD0BWP U9414 ( .A1(n3999), .A2(n3998), .ZN(n3972) );
  XNR2D1BWP U9415 ( .A1(n3951), .A2(n4712), .ZN(n3998) );
  NR2XD0BWP U9416 ( .A1(n5695), .A2(n5623), .ZN(n4712) );
  NR2XD0BWP U9417 ( .A1(n4658), .A2(n4640), .ZN(n5623) );
  NR2XD0BWP U9418 ( .A1(\alu/N684 ), .A2(\alu/N683 ), .ZN(n5695) );
  AOI21D1BWP U9419 ( .A1(op2[13]), .A2(n3653), .B(n4713), .ZN(n3951) );
  AOI21D1BWP U9420 ( .A1(n4838), .A2(n4714), .B(n4713), .ZN(n4753) );
  NR2XD0BWP U9421 ( .A1(n4714), .A2(n4838), .ZN(n4713) );
  OAI22D1BWP U9422 ( .A1(n4079), .A2(n4078), .B1(op2[12]), .B2(n4660), .ZN(
        n4714) );
  NR2XD0BWP U9423 ( .A1(n4077), .A2(op1[12]), .ZN(n4078) );
  OAI22D1BWP U9424 ( .A1(n3653), .A2(n3561), .B1(op2[13]), .B2(op1[13]), .ZN(
        n4839) );
  OR4XD1BWP U9425 ( .A1(op1[13]), .A2(\alu/N683 ), .A3(op1[12]), .A4(n5630), 
        .Z(\alu/N87 ) );
  NR2XD0BWP U9426 ( .A1(n3960), .A2(n4649), .ZN(n3952) );
  XNR3D1BWP U9427 ( .A1(op2[12]), .A2(op1[12]), .A3(n4079), .ZN(n4751) );
  AOI22D1BWP U9428 ( .A1(n5629), .A2(n3949), .B1(op1[11]), .B2(n4693), .ZN(
        n4079) );
  NR2XD0BWP U9429 ( .A1(n4676), .A2(n4677), .ZN(\intadd_36/B[0] ) );
  XOR3D1BWP U9430 ( .A1(op2[11]), .A2(n5629), .A3(n4678), .Z(n3652) );
  ND4D1BWP U9431 ( .A1(n5225), .A2(n5224), .A3(n5223), .A4(n5222), .ZN(N4205)
         );
  AOI31D1BWP U9432 ( .A1(n5217), .A2(n5219), .A3(n5218), .B(n3661), .ZN(n5220)
         );
  AOI22D1BWP U9433 ( .A1(vectorData2[157]), .A2(n5232), .B1(vectorData2[221]), 
        .B2(n5228), .ZN(n5218) );
  AOI22D1BWP U9434 ( .A1(vectorData2[173]), .A2(n5230), .B1(vectorData2[205]), 
        .B2(n5227), .ZN(n5219) );
  OA211D1BWP U9435 ( .A1(n5216), .A2(n3673), .B(n5215), .C(n5214), .Z(n5217)
         );
  AOI22D1BWP U9436 ( .A1(vectorData2[189]), .A2(n5233), .B1(vectorData2[109]), 
        .B2(n3671), .ZN(n5214) );
  AOI22D1BWP U9437 ( .A1(vectorData2[125]), .A2(n5231), .B1(vectorData2[253]), 
        .B2(n5229), .ZN(n5215) );
  AOI22D1BWP U9438 ( .A1(vectorData2[237]), .A2(n4694), .B1(scalarData2[13]), 
        .B2(n4688), .ZN(n5221) );
  INR2D1BWP U9439 ( .A1(n5187), .B1(n3661), .ZN(n4694) );
  AOI22D1BWP U9440 ( .A1(vectorData2[45]), .A2(n4687), .B1(vectorData2[93]), 
        .B2(n4684), .ZN(n5223) );
  NR2XD0BWP U9441 ( .A1(n3752), .A2(n3661), .ZN(n4684) );
  NR2XD0BWP U9442 ( .A1(n3616), .A2(n3661), .ZN(n4687) );
  AOI22D1BWP U9443 ( .A1(vectorData2[77]), .A2(n4682), .B1(vectorData2[61]), 
        .B2(n4686), .ZN(n5224) );
  NR2XD0BWP U9444 ( .A1(n3751), .A2(n3661), .ZN(n4682) );
  AOI22D1BWP U9445 ( .A1(vectorData2[29]), .A2(n4685), .B1(vectorData2[13]), 
        .B2(n4681), .ZN(n5225) );
  NR2XD0BWP U9446 ( .A1(n6063), .A2(n6043), .ZN(\vrf/N214 ) );
  NR2XD0BWP U9447 ( .A1(n6063), .A2(n6042), .ZN(\vrf/N213 ) );
  NR2XD0BWP U9448 ( .A1(n6063), .A2(n6041), .ZN(\vrf/N212 ) );
  INR2D1BWP U9449 ( .A1(vectorToLoad[192]), .B1(n6063), .ZN(\vrf/N211 ) );
  INR2D1BWP U9450 ( .A1(vectorToLoad[191]), .B1(n6063), .ZN(\vrf/N210 ) );
  INR2D1BWP U9451 ( .A1(vectorToLoad[190]), .B1(n6063), .ZN(\vrf/N209 ) );
  INR2D1BWP U9452 ( .A1(vectorToLoad[189]), .B1(n6063), .ZN(\vrf/N208 ) );
  INR2D1BWP U9453 ( .A1(vectorToLoad[188]), .B1(n6063), .ZN(\vrf/N207 ) );
  INR2D1BWP U9454 ( .A1(vectorToLoad[187]), .B1(n6063), .ZN(\vrf/N206 ) );
  INR2D1BWP U9455 ( .A1(vectorToLoad[186]), .B1(n6063), .ZN(\vrf/N205 ) );
  INR2D1BWP U9456 ( .A1(vectorToLoad[185]), .B1(n6063), .ZN(\vrf/N204 ) );
  INR2D1BWP U9457 ( .A1(vectorToLoad[184]), .B1(n6063), .ZN(\vrf/N203 ) );
  INR2D1BWP U9458 ( .A1(vectorToLoad[183]), .B1(n6063), .ZN(\vrf/N202 ) );
  INR2D1BWP U9459 ( .A1(vectorToLoad[182]), .B1(n6063), .ZN(\vrf/N201 ) );
  INR2D1BWP U9460 ( .A1(vectorToLoad[181]), .B1(n6063), .ZN(\vrf/N200 ) );
  INR2D1BWP U9461 ( .A1(vectorToLoad[180]), .B1(n6063), .ZN(\vrf/N199 ) );
  INR2D1BWP U9462 ( .A1(vectorToLoad[179]), .B1(n6063), .ZN(\vrf/N198 ) );
  INR2D1BWP U9463 ( .A1(vectorToLoad[178]), .B1(n6063), .ZN(\vrf/N197 ) );
  INR2D1BWP U9464 ( .A1(vectorToLoad[177]), .B1(n6063), .ZN(\vrf/N196 ) );
  INR2D1BWP U9465 ( .A1(vectorToLoad[176]), .B1(n6063), .ZN(\vrf/N195 ) );
  INR2D1BWP U9466 ( .A1(vectorToLoad[175]), .B1(n6063), .ZN(\vrf/N194 ) );
  INR2D1BWP U9467 ( .A1(vectorToLoad[174]), .B1(n6063), .ZN(\vrf/N193 ) );
  INR2D1BWP U9468 ( .A1(vectorToLoad[173]), .B1(n6063), .ZN(\vrf/N192 ) );
  INR2D1BWP U9469 ( .A1(vectorToLoad[172]), .B1(n6063), .ZN(\vrf/N191 ) );
  INR2D1BWP U9470 ( .A1(vectorToLoad[171]), .B1(n6063), .ZN(\vrf/N190 ) );
  INR2D1BWP U9471 ( .A1(vectorToLoad[170]), .B1(n6063), .ZN(\vrf/N189 ) );
  INR2D1BWP U9472 ( .A1(vectorToLoad[169]), .B1(n6063), .ZN(\vrf/N188 ) );
  INR2D1BWP U9473 ( .A1(vectorToLoad[168]), .B1(n6063), .ZN(\vrf/N187 ) );
  INR2D1BWP U9474 ( .A1(vectorToLoad[167]), .B1(n6063), .ZN(\vrf/N186 ) );
  INR2D1BWP U9475 ( .A1(vectorToLoad[166]), .B1(n6063), .ZN(\vrf/N185 ) );
  INR2D1BWP U9476 ( .A1(vectorToLoad[165]), .B1(n6063), .ZN(\vrf/N184 ) );
  INR2D1BWP U9477 ( .A1(vectorToLoad[164]), .B1(n6063), .ZN(\vrf/N183 ) );
  INR2D1BWP U9478 ( .A1(vectorToLoad[163]), .B1(n6063), .ZN(\vrf/N182 ) );
  INR2D1BWP U9479 ( .A1(vectorToLoad[162]), .B1(n6063), .ZN(\vrf/N181 ) );
  INR2D1BWP U9480 ( .A1(vectorToLoad[161]), .B1(n6063), .ZN(\vrf/N180 ) );
  INR2D1BWP U9481 ( .A1(vectorToLoad[160]), .B1(n6063), .ZN(\vrf/N179 ) );
  INR2D1BWP U9482 ( .A1(vectorToLoad[159]), .B1(n6063), .ZN(\vrf/N178 ) );
  INR2D1BWP U9483 ( .A1(vectorToLoad[158]), .B1(n6063), .ZN(\vrf/N177 ) );
  INR2D1BWP U9484 ( .A1(vectorToLoad[157]), .B1(n6063), .ZN(\vrf/N176 ) );
  INR2D1BWP U9485 ( .A1(vectorToLoad[156]), .B1(n6063), .ZN(\vrf/N175 ) );
  INR2D1BWP U9486 ( .A1(vectorToLoad[155]), .B1(n6063), .ZN(\vrf/N174 ) );
  INR2D1BWP U9487 ( .A1(vectorToLoad[154]), .B1(n6063), .ZN(\vrf/N173 ) );
  INR2D1BWP U9488 ( .A1(vectorToLoad[153]), .B1(n6063), .ZN(\vrf/N172 ) );
  INR2D1BWP U9489 ( .A1(vectorToLoad[152]), .B1(n6063), .ZN(\vrf/N171 ) );
  INR2D1BWP U9490 ( .A1(vectorToLoad[151]), .B1(n6063), .ZN(\vrf/N170 ) );
  INR2D1BWP U9491 ( .A1(vectorToLoad[150]), .B1(n6063), .ZN(\vrf/N169 ) );
  INR2D1BWP U9492 ( .A1(vectorToLoad[149]), .B1(n6063), .ZN(\vrf/N168 ) );
  INR2D1BWP U9493 ( .A1(vectorToLoad[148]), .B1(n6063), .ZN(\vrf/N167 ) );
  INR2D1BWP U9494 ( .A1(vectorToLoad[147]), .B1(n6063), .ZN(\vrf/N166 ) );
  NR2XD0BWP U9495 ( .A1(n4997), .A2(n4993), .ZN(n5185) );
  ND3D1BWP U9496 ( .A1(n4698), .A2(n3679), .A3(n5417), .ZN(n4997) );
  ND3D1BWP U9497 ( .A1(cycles[1]), .A2(n4698), .A3(n3679), .ZN(n4995) );
  NR2XD0BWP U9498 ( .A1(n4999), .A2(n4993), .ZN(n5213) );
  ND3D1BWP U9499 ( .A1(cycles[0]), .A2(n4698), .A3(n5417), .ZN(n4999) );
  NR2XD0BWP U9500 ( .A1(n3748), .A2(n3749), .ZN(n4681) );
  AOI21D1BWP U9501 ( .A1(n3746), .A2(n3745), .B(n3944), .ZN(n3883) );
  INR2D1BWP U9502 ( .A1(n3787), .B1(n3749), .ZN(n3944) );
  INR2D1BWP U9503 ( .A1(vectorToLoad[41]), .B1(n6063), .ZN(\vrf/N59 ) );
  INR2D1BWP U9504 ( .A1(vectorToLoad[40]), .B1(n6063), .ZN(\vrf/N58 ) );
  INR2D1BWP U9505 ( .A1(vectorToLoad[39]), .B1(n6063), .ZN(\vrf/N57 ) );
  INR2D1BWP U9506 ( .A1(vectorToLoad[38]), .B1(n6063), .ZN(\vrf/N56 ) );
  INR2D1BWP U9507 ( .A1(vectorToLoad[37]), .B1(n6063), .ZN(\vrf/N55 ) );
  INR2D1BWP U9508 ( .A1(vectorToLoad[36]), .B1(n6063), .ZN(\vrf/N54 ) );
  INR2D1BWP U9509 ( .A1(vectorToLoad[35]), .B1(n6063), .ZN(\vrf/N53 ) );
  INR2D1BWP U9510 ( .A1(vectorToLoad[34]), .B1(n6063), .ZN(\vrf/N52 ) );
  INR2D1BWP U9511 ( .A1(vectorToLoad[33]), .B1(n6063), .ZN(\vrf/N51 ) );
  INR2D1BWP U9512 ( .A1(vectorToLoad[32]), .B1(n6063), .ZN(\vrf/N50 ) );
  INR2D1BWP U9513 ( .A1(vectorToLoad[31]), .B1(n6063), .ZN(\vrf/N49 ) );
  INR2D1BWP U9514 ( .A1(vectorToLoad[30]), .B1(n6063), .ZN(\vrf/N48 ) );
  INR2D1BWP U9515 ( .A1(vectorToLoad[29]), .B1(n6063), .ZN(\vrf/N47 ) );
  INR2D1BWP U9516 ( .A1(vectorToLoad[28]), .B1(n6063), .ZN(\vrf/N46 ) );
  INR2D1BWP U9517 ( .A1(vectorToLoad[27]), .B1(n6063), .ZN(\vrf/N45 ) );
  INR2D1BWP U9518 ( .A1(vectorToLoad[26]), .B1(n6063), .ZN(\vrf/N44 ) );
  INR2D1BWP U9519 ( .A1(vectorToLoad[25]), .B1(n6063), .ZN(\vrf/N43 ) );
  INR2D1BWP U9520 ( .A1(vectorToLoad[24]), .B1(n6063), .ZN(\vrf/N42 ) );
  INR2D1BWP U9521 ( .A1(vectorToLoad[23]), .B1(n6063), .ZN(\vrf/N41 ) );
  INR2D1BWP U9522 ( .A1(vectorToLoad[22]), .B1(n6063), .ZN(\vrf/N40 ) );
  INR2D1BWP U9523 ( .A1(vectorToLoad[21]), .B1(n6063), .ZN(\vrf/N39 ) );
  INR2D1BWP U9524 ( .A1(vectorToLoad[20]), .B1(n6063), .ZN(\vrf/N38 ) );
  INR2D1BWP U9525 ( .A1(vectorToLoad[19]), .B1(n6063), .ZN(\vrf/N37 ) );
  INR2D1BWP U9526 ( .A1(vectorToLoad[18]), .B1(n6063), .ZN(\vrf/N36 ) );
  INR2D1BWP U9527 ( .A1(vectorToLoad[17]), .B1(n6063), .ZN(\vrf/N35 ) );
  INR2D1BWP U9528 ( .A1(vectorToLoad[16]), .B1(n6063), .ZN(\vrf/N34 ) );
  NR2XD0BWP U9529 ( .A1(n6063), .A2(n113), .ZN(\vrf/N33 ) );
  NR2XD0BWP U9530 ( .A1(n6063), .A2(n114), .ZN(\vrf/N32 ) );
  NR2XD0BWP U9531 ( .A1(n6063), .A2(n115), .ZN(\vrf/N31 ) );
  NR2XD0BWP U9532 ( .A1(n6063), .A2(n116), .ZN(\vrf/N30 ) );
  NR2XD0BWP U9533 ( .A1(n6063), .A2(n117), .ZN(\vrf/N29 ) );
  NR2XD0BWP U9534 ( .A1(n6063), .A2(n118), .ZN(\vrf/N28 ) );
  NR2XD0BWP U9535 ( .A1(n6063), .A2(n119), .ZN(\vrf/N27 ) );
  NR2XD0BWP U9536 ( .A1(n6063), .A2(n120), .ZN(\vrf/N26 ) );
  NR2XD0BWP U9537 ( .A1(n6063), .A2(n121), .ZN(\vrf/N25 ) );
  NR2XD0BWP U9538 ( .A1(n6063), .A2(n122), .ZN(\vrf/N24 ) );
  NR2XD0BWP U9539 ( .A1(n6063), .A2(n123), .ZN(\vrf/N23 ) );
  NR2XD0BWP U9540 ( .A1(n6063), .A2(n124), .ZN(\vrf/N22 ) );
  NR2XD0BWP U9541 ( .A1(n6063), .A2(n125), .ZN(\vrf/N21 ) );
  NR2XD0BWP U9542 ( .A1(n6063), .A2(n126), .ZN(\vrf/N20 ) );
  NR2XD0BWP U9543 ( .A1(n6063), .A2(n127), .ZN(\vrf/N19 ) );
  NR2XD0BWP U9544 ( .A1(n6063), .A2(n128), .ZN(\vrf/N18 ) );
  INR2D1BWP U9545 ( .A1(vectorToLoad[255]), .B1(n6063), .ZN(\vrf/N275 ) );
  INR2D1BWP U9546 ( .A1(vectorToLoad[254]), .B1(n6063), .ZN(\vrf/N274 ) );
  INR2D1BWP U9547 ( .A1(vectorToLoad[253]), .B1(n6063), .ZN(\vrf/N273 ) );
  INR2D1BWP U9548 ( .A1(vectorToLoad[252]), .B1(n6063), .ZN(\vrf/N272 ) );
  INR2D1BWP U9549 ( .A1(vectorToLoad[251]), .B1(n6063), .ZN(\vrf/N271 ) );
  INR2D1BWP U9550 ( .A1(vectorToLoad[250]), .B1(n6063), .ZN(\vrf/N270 ) );
  INR2D1BWP U9551 ( .A1(vectorToLoad[249]), .B1(n6063), .ZN(\vrf/N269 ) );
  INR2D1BWP U9552 ( .A1(vectorToLoad[248]), .B1(n6063), .ZN(\vrf/N268 ) );
  INR2D1BWP U9553 ( .A1(vectorToLoad[247]), .B1(n6063), .ZN(\vrf/N267 ) );
  INR2D1BWP U9554 ( .A1(vectorToLoad[42]), .B1(n6063), .ZN(\vrf/N60 ) );
  INR2D1BWP U9555 ( .A1(vectorToLoad[246]), .B1(n6063), .ZN(\vrf/N266 ) );
  INR2D1BWP U9556 ( .A1(vectorToLoad[245]), .B1(n6063), .ZN(\vrf/N265 ) );
  INR2D1BWP U9557 ( .A1(vectorToLoad[244]), .B1(n6063), .ZN(\vrf/N264 ) );
  INR2D1BWP U9558 ( .A1(vectorToLoad[243]), .B1(n6063), .ZN(\vrf/N263 ) );
  INR2D1BWP U9559 ( .A1(vectorToLoad[242]), .B1(n6063), .ZN(\vrf/N262 ) );
  INR2D1BWP U9560 ( .A1(vectorToLoad[241]), .B1(n6063), .ZN(\vrf/N261 ) );
  INR2D1BWP U9561 ( .A1(vectorToLoad[240]), .B1(n6063), .ZN(\vrf/N260 ) );
  INR2D1BWP U9562 ( .A1(vectorToLoad[239]), .B1(n6063), .ZN(\vrf/N259 ) );
  INR2D1BWP U9563 ( .A1(vectorToLoad[238]), .B1(n6063), .ZN(\vrf/N258 ) );
  INR2D1BWP U9564 ( .A1(vectorToLoad[237]), .B1(n6063), .ZN(\vrf/N257 ) );
  INR2D1BWP U9565 ( .A1(vectorToLoad[236]), .B1(n6063), .ZN(\vrf/N256 ) );
  INR2D1BWP U9566 ( .A1(vectorToLoad[235]), .B1(n6063), .ZN(\vrf/N255 ) );
  INR2D1BWP U9567 ( .A1(vectorToLoad[234]), .B1(n6063), .ZN(\vrf/N254 ) );
  INR2D1BWP U9568 ( .A1(vectorToLoad[233]), .B1(n6063), .ZN(\vrf/N253 ) );
  INR2D1BWP U9569 ( .A1(vectorToLoad[232]), .B1(n6063), .ZN(\vrf/N252 ) );
  INR2D1BWP U9570 ( .A1(vectorToLoad[231]), .B1(n6063), .ZN(\vrf/N251 ) );
  INR2D1BWP U9571 ( .A1(vectorToLoad[230]), .B1(n6063), .ZN(\vrf/N250 ) );
  INR2D1BWP U9572 ( .A1(vectorToLoad[229]), .B1(n6063), .ZN(\vrf/N249 ) );
  INR2D1BWP U9573 ( .A1(vectorToLoad[228]), .B1(n6063), .ZN(\vrf/N248 ) );
  INR2D1BWP U9574 ( .A1(vectorToLoad[227]), .B1(n6063), .ZN(\vrf/N247 ) );
  INR2D1BWP U9575 ( .A1(vectorToLoad[226]), .B1(n6063), .ZN(\vrf/N246 ) );
  INR2D1BWP U9576 ( .A1(vectorToLoad[225]), .B1(n6063), .ZN(\vrf/N245 ) );
  INR2D1BWP U9577 ( .A1(vectorToLoad[224]), .B1(n6063), .ZN(\vrf/N244 ) );
  NR2XD0BWP U9578 ( .A1(n6063), .A2(n6061), .ZN(\vrf/N243 ) );
  NR2XD0BWP U9579 ( .A1(n6063), .A2(n6060), .ZN(\vrf/N242 ) );
  INR2D1BWP U9580 ( .A1(vectorToLoad[221]), .B1(n6063), .ZN(\vrf/N241 ) );
  NR2XD0BWP U9581 ( .A1(n6063), .A2(n6059), .ZN(\vrf/N240 ) );
  NR2XD0BWP U9582 ( .A1(n6063), .A2(n6058), .ZN(\vrf/N239 ) );
  NR2XD0BWP U9583 ( .A1(n6063), .A2(n6057), .ZN(\vrf/N238 ) );
  NR2XD0BWP U9584 ( .A1(n6063), .A2(n6056), .ZN(\vrf/N237 ) );
  NR2XD0BWP U9585 ( .A1(n6063), .A2(n6055), .ZN(\vrf/N236 ) );
  NR2XD0BWP U9586 ( .A1(n6063), .A2(n6054), .ZN(\vrf/N235 ) );
  NR2XD0BWP U9587 ( .A1(n6063), .A2(n6053), .ZN(\vrf/N234 ) );
  INR2D1BWP U9588 ( .A1(vectorToLoad[213]), .B1(n6063), .ZN(\vrf/N233 ) );
  NR2XD0BWP U9589 ( .A1(n6063), .A2(n6052), .ZN(\vrf/N232 ) );
  NR2XD0BWP U9590 ( .A1(n6063), .A2(n6051), .ZN(\vrf/N231 ) );
  INR2D1BWP U9591 ( .A1(vectorToLoad[210]), .B1(n6063), .ZN(\vrf/N230 ) );
  NR2XD0BWP U9592 ( .A1(n6063), .A2(n6050), .ZN(\vrf/N229 ) );
  INR2D1BWP U9593 ( .A1(vectorToLoad[208]), .B1(n6063), .ZN(\vrf/N228 ) );
  NR2XD0BWP U9594 ( .A1(n6063), .A2(n6049), .ZN(\vrf/N227 ) );
  INR2D1BWP U9595 ( .A1(vectorToLoad[206]), .B1(n6063), .ZN(\vrf/N226 ) );
  NR2XD0BWP U9596 ( .A1(n6063), .A2(n6048), .ZN(\vrf/N225 ) );
  NR2XD0BWP U9597 ( .A1(n6063), .A2(n6047), .ZN(\vrf/N224 ) );
  NR2XD0BWP U9598 ( .A1(n6063), .A2(n6046), .ZN(\vrf/N223 ) );
  INR2D1BWP U9599 ( .A1(vectorToLoad[202]), .B1(n6063), .ZN(\vrf/N222 ) );
  NR2XD0BWP U9600 ( .A1(n6063), .A2(n6045), .ZN(\vrf/N221 ) );
  INR2D1BWP U9601 ( .A1(vectorToLoad[200]), .B1(n6063), .ZN(\vrf/N220 ) );
  INR2D1BWP U9602 ( .A1(vectorToLoad[199]), .B1(n6063), .ZN(\vrf/N219 ) );
  INR2D1BWP U9603 ( .A1(vectorToLoad[198]), .B1(n6063), .ZN(\vrf/N218 ) );
  NR2XD0BWP U9604 ( .A1(n6063), .A2(n6044), .ZN(\vrf/N216 ) );
  INR2D1BWP U9605 ( .A1(vectorToLoad[196]), .B1(n6063), .ZN(\vrf/N215 ) );
  INR2D1BWP U9606 ( .A1(vectorToLoad[43]), .B1(n6063), .ZN(\vrf/N61 ) );
  INR2D1BWP U9607 ( .A1(vectorToLoad[145]), .B1(n6063), .ZN(\vrf/N164 ) );
  INR2D1BWP U9608 ( .A1(vectorToLoad[144]), .B1(n6063), .ZN(\vrf/N163 ) );
  INR2D1BWP U9609 ( .A1(vectorToLoad[143]), .B1(n6063), .ZN(\vrf/N162 ) );
  INR2D1BWP U9610 ( .A1(vectorToLoad[142]), .B1(n6063), .ZN(\vrf/N161 ) );
  INR2D1BWP U9611 ( .A1(vectorToLoad[141]), .B1(n6063), .ZN(\vrf/N160 ) );
  INR2D1BWP U9612 ( .A1(vectorToLoad[140]), .B1(n6063), .ZN(\vrf/N159 ) );
  INR2D1BWP U9613 ( .A1(vectorToLoad[139]), .B1(n6063), .ZN(\vrf/N158 ) );
  INR2D1BWP U9614 ( .A1(vectorToLoad[138]), .B1(n6063), .ZN(\vrf/N157 ) );
  INR2D1BWP U9615 ( .A1(vectorToLoad[137]), .B1(n6063), .ZN(\vrf/N156 ) );
  INR2D1BWP U9616 ( .A1(vectorToLoad[136]), .B1(n6063), .ZN(\vrf/N155 ) );
  INR2D1BWP U9617 ( .A1(vectorToLoad[135]), .B1(n6063), .ZN(\vrf/N154 ) );
  INR2D1BWP U9618 ( .A1(vectorToLoad[134]), .B1(n6063), .ZN(\vrf/N153 ) );
  INR2D1BWP U9619 ( .A1(vectorToLoad[133]), .B1(n6063), .ZN(\vrf/N152 ) );
  INR2D1BWP U9620 ( .A1(vectorToLoad[132]), .B1(n6063), .ZN(\vrf/N151 ) );
  INR2D1BWP U9621 ( .A1(vectorToLoad[131]), .B1(n6063), .ZN(\vrf/N150 ) );
  INR2D1BWP U9622 ( .A1(vectorToLoad[130]), .B1(n6063), .ZN(\vrf/N149 ) );
  INR2D1BWP U9623 ( .A1(vectorToLoad[129]), .B1(n6063), .ZN(\vrf/N148 ) );
  INR2D1BWP U9624 ( .A1(vectorToLoad[128]), .B1(n6063), .ZN(\vrf/N147 ) );
  INR2D1BWP U9625 ( .A1(vectorToLoad[127]), .B1(n6063), .ZN(\vrf/N146 ) );
  INR2D1BWP U9626 ( .A1(vectorToLoad[126]), .B1(n6063), .ZN(\vrf/N145 ) );
  INR2D1BWP U9627 ( .A1(vectorToLoad[125]), .B1(n6063), .ZN(\vrf/N144 ) );
  INR2D1BWP U9628 ( .A1(vectorToLoad[124]), .B1(n6063), .ZN(\vrf/N143 ) );
  INR2D1BWP U9629 ( .A1(vectorToLoad[123]), .B1(n6063), .ZN(\vrf/N142 ) );
  INR2D1BWP U9630 ( .A1(vectorToLoad[122]), .B1(n6063), .ZN(\vrf/N141 ) );
  INR2D1BWP U9631 ( .A1(vectorToLoad[121]), .B1(n6063), .ZN(\vrf/N140 ) );
  INR2D1BWP U9632 ( .A1(vectorToLoad[120]), .B1(n6063), .ZN(\vrf/N139 ) );
  INR2D1BWP U9633 ( .A1(vectorToLoad[119]), .B1(n6063), .ZN(\vrf/N138 ) );
  INR2D1BWP U9634 ( .A1(vectorToLoad[118]), .B1(n6063), .ZN(\vrf/N137 ) );
  INR2D1BWP U9635 ( .A1(vectorToLoad[117]), .B1(n6063), .ZN(\vrf/N136 ) );
  INR2D1BWP U9636 ( .A1(vectorToLoad[116]), .B1(n6063), .ZN(\vrf/N135 ) );
  INR2D1BWP U9637 ( .A1(vectorToLoad[115]), .B1(n6063), .ZN(\vrf/N134 ) );
  INR2D1BWP U9638 ( .A1(vectorToLoad[114]), .B1(n6063), .ZN(\vrf/N133 ) );
  INR2D1BWP U9639 ( .A1(vectorToLoad[113]), .B1(n6063), .ZN(\vrf/N132 ) );
  INR2D1BWP U9640 ( .A1(vectorToLoad[112]), .B1(n6063), .ZN(\vrf/N131 ) );
  INR2D1BWP U9641 ( .A1(vectorToLoad[111]), .B1(n6063), .ZN(\vrf/N130 ) );
  INR2D1BWP U9642 ( .A1(vectorToLoad[110]), .B1(n6063), .ZN(\vrf/N129 ) );
  INR2D1BWP U9643 ( .A1(vectorToLoad[109]), .B1(n6063), .ZN(\vrf/N128 ) );
  INR2D1BWP U9644 ( .A1(vectorToLoad[108]), .B1(n6063), .ZN(\vrf/N127 ) );
  INR2D1BWP U9645 ( .A1(vectorToLoad[107]), .B1(n6063), .ZN(\vrf/N126 ) );
  INR2D1BWP U9646 ( .A1(vectorToLoad[106]), .B1(n6063), .ZN(\vrf/N125 ) );
  INR2D1BWP U9647 ( .A1(vectorToLoad[105]), .B1(n6063), .ZN(\vrf/N124 ) );
  INR2D1BWP U9648 ( .A1(vectorToLoad[104]), .B1(n6063), .ZN(\vrf/N123 ) );
  INR2D1BWP U9649 ( .A1(vectorToLoad[103]), .B1(n6063), .ZN(\vrf/N122 ) );
  INR2D1BWP U9650 ( .A1(vectorToLoad[102]), .B1(n6063), .ZN(\vrf/N121 ) );
  INR2D1BWP U9651 ( .A1(vectorToLoad[101]), .B1(n6063), .ZN(\vrf/N120 ) );
  INR2D1BWP U9652 ( .A1(vectorToLoad[100]), .B1(n6063), .ZN(\vrf/N119 ) );
  INR2D1BWP U9653 ( .A1(vectorToLoad[99]), .B1(n6063), .ZN(\vrf/N118 ) );
  INR2D1BWP U9654 ( .A1(vectorToLoad[98]), .B1(n6063), .ZN(\vrf/N116 ) );
  INR2D1BWP U9655 ( .A1(vectorToLoad[97]), .B1(n6063), .ZN(\vrf/N115 ) );
  INR2D1BWP U9656 ( .A1(vectorToLoad[96]), .B1(n6063), .ZN(\vrf/N114 ) );
  INR2D1BWP U9657 ( .A1(vectorToLoad[95]), .B1(n6063), .ZN(\vrf/N113 ) );
  INR2D1BWP U9658 ( .A1(vectorToLoad[94]), .B1(n6063), .ZN(\vrf/N112 ) );
  INR2D1BWP U9659 ( .A1(vectorToLoad[44]), .B1(n6063), .ZN(\vrf/N62 ) );
  INR2D1BWP U9660 ( .A1(vectorToLoad[45]), .B1(n6063), .ZN(\vrf/N63 ) );
  INR2D1BWP U9661 ( .A1(vectorToLoad[46]), .B1(n6063), .ZN(\vrf/N64 ) );
  INR2D1BWP U9662 ( .A1(vectorToLoad[47]), .B1(n6063), .ZN(\vrf/N65 ) );
  INR2D1BWP U9663 ( .A1(vectorToLoad[48]), .B1(n6063), .ZN(\vrf/N66 ) );
  INR2D1BWP U9664 ( .A1(vectorToLoad[49]), .B1(n6063), .ZN(\vrf/N67 ) );
  INR2D1BWP U9665 ( .A1(vectorToLoad[50]), .B1(n6063), .ZN(\vrf/N68 ) );
  INR2D1BWP U9666 ( .A1(vectorToLoad[51]), .B1(n6063), .ZN(\vrf/N69 ) );
  INR2D1BWP U9667 ( .A1(vectorToLoad[52]), .B1(n6063), .ZN(\vrf/N70 ) );
  INR2D1BWP U9668 ( .A1(vectorToLoad[53]), .B1(n6063), .ZN(\vrf/N71 ) );
  INR2D1BWP U9669 ( .A1(vectorToLoad[54]), .B1(n6063), .ZN(\vrf/N72 ) );
  INR2D1BWP U9670 ( .A1(vectorToLoad[55]), .B1(n6063), .ZN(\vrf/N73 ) );
  INR2D1BWP U9671 ( .A1(vectorToLoad[57]), .B1(n6063), .ZN(\vrf/N75 ) );
  INR2D1BWP U9672 ( .A1(vectorToLoad[58]), .B1(n6063), .ZN(\vrf/N76 ) );
  INR2D1BWP U9673 ( .A1(vectorToLoad[59]), .B1(n6063), .ZN(\vrf/N77 ) );
  INR2D1BWP U9674 ( .A1(vectorToLoad[60]), .B1(n6063), .ZN(\vrf/N78 ) );
  INR2D1BWP U9675 ( .A1(vectorToLoad[61]), .B1(n6063), .ZN(\vrf/N79 ) );
  INR2D1BWP U9676 ( .A1(vectorToLoad[62]), .B1(n6063), .ZN(\vrf/N80 ) );
  INR2D1BWP U9677 ( .A1(vectorToLoad[63]), .B1(n6063), .ZN(\vrf/N81 ) );
  INR2D1BWP U9678 ( .A1(vectorToLoad[64]), .B1(n6063), .ZN(\vrf/N82 ) );
  INR2D1BWP U9679 ( .A1(vectorToLoad[65]), .B1(n6063), .ZN(\vrf/N83 ) );
  INR2D1BWP U9680 ( .A1(vectorToLoad[66]), .B1(n6063), .ZN(\vrf/N84 ) );
  INR2D1BWP U9681 ( .A1(vectorToLoad[67]), .B1(n6063), .ZN(\vrf/N85 ) );
  INR2D1BWP U9682 ( .A1(vectorToLoad[68]), .B1(n6063), .ZN(\vrf/N86 ) );
  INR2D1BWP U9683 ( .A1(vectorToLoad[69]), .B1(n6063), .ZN(\vrf/N87 ) );
  INR2D1BWP U9684 ( .A1(vectorToLoad[70]), .B1(n6063), .ZN(\vrf/N88 ) );
  INR2D1BWP U9685 ( .A1(vectorToLoad[71]), .B1(n6063), .ZN(\vrf/N89 ) );
  INR2D1BWP U9686 ( .A1(vectorToLoad[72]), .B1(n6063), .ZN(\vrf/N90 ) );
  INR2D1BWP U9687 ( .A1(vectorToLoad[73]), .B1(n6063), .ZN(\vrf/N91 ) );
  INR2D1BWP U9688 ( .A1(vectorToLoad[74]), .B1(n6063), .ZN(\vrf/N92 ) );
  INR2D1BWP U9689 ( .A1(vectorToLoad[75]), .B1(n6063), .ZN(\vrf/N93 ) );
  INR2D1BWP U9690 ( .A1(vectorToLoad[76]), .B1(n6063), .ZN(\vrf/N94 ) );
  INR2D1BWP U9691 ( .A1(vectorToLoad[77]), .B1(n6063), .ZN(\vrf/N95 ) );
  INR2D1BWP U9692 ( .A1(vectorToLoad[78]), .B1(n6063), .ZN(\vrf/N96 ) );
  INR2D1BWP U9693 ( .A1(vectorToLoad[79]), .B1(n6063), .ZN(\vrf/N97 ) );
  INR2D1BWP U9694 ( .A1(vectorToLoad[80]), .B1(n6063), .ZN(\vrf/N98 ) );
  INR2D1BWP U9695 ( .A1(vectorToLoad[81]), .B1(n6063), .ZN(\vrf/N99 ) );
  INR2D1BWP U9696 ( .A1(vectorToLoad[146]), .B1(n6063), .ZN(\vrf/N165 ) );
  INR2D1BWP U9697 ( .A1(vectorToLoad[56]), .B1(n6063), .ZN(\vrf/N74 ) );
  INR2D1BWP U9698 ( .A1(vectorToLoad[91]), .B1(n6063), .ZN(\vrf/N109 ) );
  INR2D1BWP U9699 ( .A1(vectorToLoad[82]), .B1(n6063), .ZN(\vrf/N100 ) );
  INR2D1BWP U9700 ( .A1(vectorToLoad[83]), .B1(n6063), .ZN(\vrf/N101 ) );
  INR2D1BWP U9701 ( .A1(vectorToLoad[85]), .B1(n6063), .ZN(\vrf/N103 ) );
  INR2D1BWP U9702 ( .A1(vectorToLoad[87]), .B1(n6063), .ZN(\vrf/N105 ) );
  INR2D1BWP U9703 ( .A1(vectorToLoad[88]), .B1(n6063), .ZN(\vrf/N106 ) );
  INR2D1BWP U9704 ( .A1(vectorToLoad[92]), .B1(n6063), .ZN(\vrf/N110 ) );
  INR2D1BWP U9705 ( .A1(vectorToLoad[90]), .B1(n6063), .ZN(\vrf/N108 ) );
  INR2D1BWP U9706 ( .A1(vectorToLoad[89]), .B1(n6063), .ZN(\vrf/N107 ) );
  INR2D1BWP U9707 ( .A1(vectorToLoad[86]), .B1(n6063), .ZN(\vrf/N104 ) );
  INR2D1BWP U9708 ( .A1(vectorToLoad[84]), .B1(n6063), .ZN(\vrf/N102 ) );
  INR2D1BWP U9709 ( .A1(vectorToLoad[93]), .B1(n6063), .ZN(\vrf/N111 ) );
  NR2XD0BWP U9710 ( .A1(n5559), .A2(n5560), .ZN(\mult_x_153/n105 ) );
  AOI22D1BWP U9711 ( .A1(n4815), .A2(n4818), .B1(n4787), .B2(n4820), .ZN(n5560) );
  OAI32D1BWP U9712 ( .A1(op2[0]), .A2(op1[4]), .A3(n4832), .B1(n4680), .B2(
        n4809), .ZN(n4787) );
  IND2D1BWP U9713 ( .A1(\mult_x_153/n149 ), .B1(n5587), .ZN(n5559) );
  OAI22D1BWP U9714 ( .A1(n4792), .A2(n4793), .B1(n5554), .B2(n4791), .ZN(
        \mult_x_153/n130 ) );
  OAI22D1BWP U9715 ( .A1(n4820), .A2(n4812), .B1(n4816), .B2(n4813), .ZN(
        \mult_x_153/n154 ) );
  OAI22D1BWP U9716 ( .A1(n4792), .A2(n5554), .B1(n4793), .B2(n4794), .ZN(
        \mult_x_153/n131 ) );
  AOI22D1BWP U9717 ( .A1(op1[9]), .A2(n5569), .B1(op2[3]), .B2(n3680), .ZN(
        n4794) );
  AOI22D1BWP U9718 ( .A1(op1[9]), .A2(n4667), .B1(op2[4]), .B2(n3680), .ZN(
        n4792) );
  OAI22D1BWP U9719 ( .A1(op1[9]), .A2(n5554), .B1(n4845), .B2(n4793), .ZN(
        \mult_x_153/n125 ) );
  OAI21D1BWP U9720 ( .A1(n4662), .A2(n4832), .B(op1[7]), .ZN(\mult_x_153/n136 ) );
  AOI22D1BWP U9721 ( .A1(n4800), .A2(n4785), .B1(n4784), .B2(n4808), .ZN(n4786) );
  OAI32D1BWP U9722 ( .A1(op2[0]), .A2(op1[6]), .A3(n5605), .B1(n4680), .B2(
        n4798), .ZN(n4784) );
  AOI22D1BWP U9723 ( .A1(n5555), .A2(n4788), .B1(n4796), .B2(n4790), .ZN(n4764) );
  AOI22D1BWP U9724 ( .A1(n4800), .A2(n4762), .B1(n4806), .B2(n4799), .ZN(n4765) );
  OAI22D1BWP U9725 ( .A1(n5576), .A2(n4825), .B1(n4826), .B2(n5562), .ZN(
        \mult_x_153/n169 ) );
  AOI22D1BWP U9726 ( .A1(op1[3]), .A2(n4667), .B1(op2[4]), .B2(n5561), .ZN(
        n4826) );
  OAI22D1BWP U9727 ( .A1(n4789), .A2(n4793), .B1(n5554), .B2(n4845), .ZN(
        \mult_x_153/n126 ) );
  OAI22D1BWP U9728 ( .A1(n3680), .A2(op2[9]), .B1(n4648), .B2(op1[9]), .ZN(
        n4844) );
  OAI21D1BWP U9729 ( .A1(op2[9]), .A2(n5564), .B(n4827), .ZN(\mult_x_153/n177 ) );
  AOI22D1BWP U9730 ( .A1(n4762), .A2(n4806), .B1(n4800), .B2(n5605), .ZN(n4758) );
  AOI22D1BWP U9731 ( .A1(op1[7]), .A2(op2[9]), .B1(n4648), .B2(n5605), .ZN(
        n4762) );
  AOI22D1BWP U9732 ( .A1(op1[9]), .A2(op2[5]), .B1(op2[6]), .B2(n3680), .ZN(
        n4759) );
  OAI22D1BWP U9733 ( .A1(n3680), .A2(n4667), .B1(n5615), .B2(op1[9]), .ZN(
        n4766) );
  OAI22D1BWP U9734 ( .A1(op1[5]), .A2(n4820), .B1(n4810), .B2(n4816), .ZN(
        \mult_x_153/n151 ) );
  AOI22D1BWP U9735 ( .A1(op1[5]), .A2(n4648), .B1(op2[9]), .B2(n4832), .ZN(
        n4810) );
  AOI22D1BWP U9736 ( .A1(op1[5]), .A2(op2[1]), .B1(n5616), .B2(n4832), .ZN(
        n4818) );
  AOI22D1BWP U9737 ( .A1(n4800), .A2(n4805), .B1(n4806), .B2(n4777), .ZN(n4770) );
  AOI22D1BWP U9738 ( .A1(n4824), .A2(n5557), .B1(n4822), .B2(n5572), .ZN(n4771) );
  AOI22D1BWP U9739 ( .A1(n4815), .A2(n4852), .B1(n4817), .B2(n4778), .ZN(n4772) );
  OAI32D1BWP U9740 ( .A1(op1[3]), .A2(n6070), .A3(n4669), .B1(n5576), .B2(
        n5561), .ZN(\mult_x_153/n163 ) );
  AOI22D1BWP U9741 ( .A1(n4815), .A2(n4778), .B1(n4817), .B2(n4814), .ZN(n4780) );
  AOI22D1BWP U9742 ( .A1(op1[5]), .A2(op2[4]), .B1(n4667), .B2(n4832), .ZN(
        n4778) );
  AOI22D1BWP U9743 ( .A1(n4800), .A2(n4777), .B1(n4785), .B2(n4806), .ZN(n4781) );
  AOI22D1BWP U9744 ( .A1(op1[7]), .A2(op2[1]), .B1(n5616), .B2(n5605), .ZN(
        n4785) );
  AOI22D1BWP U9745 ( .A1(op1[7]), .A2(op2[2]), .B1(n4670), .B2(n5605), .ZN(
        n4777) );
  NR2XD0BWP U9746 ( .A1(n4808), .A2(n4680), .ZN(\mult_x_153/n148 ) );
  OAI22D1BWP U9747 ( .A1(n4808), .A2(n4801), .B1(n4803), .B2(n4802), .ZN(
        \mult_x_153/n141 ) );
  AOI22D1BWP U9748 ( .A1(op1[9]), .A2(n4680), .B1(n5616), .B2(n3680), .ZN(
        \mult_x_153/n121 ) );
  AOI22D1BWP U9749 ( .A1(n4815), .A2(n4832), .B1(n4809), .B2(n4820), .ZN(
        \mult_x_153/n150 ) );
  AOI22D1BWP U9750 ( .A1(op1[9]), .A2(n4670), .B1(n5569), .B2(n3680), .ZN(
        \mult_x_153/n120 ) );
  AOI22D1BWP U9751 ( .A1(op1[7]), .A2(op2[8]), .B1(n4654), .B2(n5605), .ZN(
        n4799) );
  OAI22D1BWP U9752 ( .A1(n5605), .A2(op2[7]), .B1(n4833), .B2(op1[7]), .ZN(
        n4849) );
  OAI21D1BWP U9753 ( .A1(op2[6]), .A2(n5564), .B(n4830), .ZN(\mult_x_153/n180 ) );
  AOI22D1BWP U9754 ( .A1(op2[7]), .A2(n5570), .B1(\mult_x_153/n176 ), .B2(
        n4833), .ZN(n4830) );
  OAI22D1BWP U9755 ( .A1(n5576), .A2(n4821), .B1(n4823), .B2(n5562), .ZN(
        \mult_x_153/n165 ) );
  OAI21D1BWP U9756 ( .A1(op2[8]), .A2(n5564), .B(n4828), .ZN(\mult_x_153/n178 ) );
  AOI22D1BWP U9757 ( .A1(op2[9]), .A2(n5570), .B1(\mult_x_153/n176 ), .B2(
        n4648), .ZN(n4828) );
  AOI22D1BWP U9758 ( .A1(op1[3]), .A2(op2[7]), .B1(n4833), .B2(n5561), .ZN(
        n4822) );
  AOI22D1BWP U9759 ( .A1(op1[3]), .A2(n4654), .B1(op2[8]), .B2(n5561), .ZN(
        n4823) );
  AOI22D1BWP U9760 ( .A1(op1[9]), .A2(op2[7]), .B1(n4833), .B2(n3680), .ZN(
        n4788) );
  AOI22D1BWP U9761 ( .A1(op1[9]), .A2(n4654), .B1(op2[8]), .B2(n3680), .ZN(
        n4789) );
  OAI21D1BWP U9762 ( .A1(op2[7]), .A2(n5564), .B(n4829), .ZN(\mult_x_153/n179 ) );
  AOI22D1BWP U9763 ( .A1(op2[8]), .A2(n5570), .B1(\mult_x_153/n176 ), .B2(
        n4654), .ZN(n4829) );
  OAI22D1BWP U9764 ( .A1(op1[3]), .A2(n5576), .B1(n4821), .B2(n5562), .ZN(
        \mult_x_153/n164 ) );
  AOI22D1BWP U9765 ( .A1(op1[3]), .A2(n4648), .B1(op2[9]), .B2(n5561), .ZN(
        n4821) );
  OAI22D1BWP U9766 ( .A1(n3680), .A2(n4663), .B1(n4833), .B2(op1[9]), .ZN(
        n6072) );
  OAI22D1BWP U9767 ( .A1(n4820), .A2(n4811), .B1(n4816), .B2(n4812), .ZN(
        \mult_x_153/n153 ) );
  AOI22D1BWP U9768 ( .A1(op1[5]), .A2(n4833), .B1(op2[7]), .B2(n4832), .ZN(
        n4812) );
  AOI22D1BWP U9769 ( .A1(op1[5]), .A2(n4654), .B1(op2[8]), .B2(n4832), .ZN(
        n4811) );
  OAI21D1BWP U9770 ( .A1(n4666), .A2(n5561), .B(op1[5]), .ZN(\mult_x_153/n149 ) );
  AOI22D1BWP U9771 ( .A1(op1[5]), .A2(op2[3]), .B1(n5569), .B2(n4832), .ZN(
        n4814) );
  AOI22D1BWP U9772 ( .A1(op1[5]), .A2(n4670), .B1(op2[2]), .B2(n4832), .ZN(
        n4819) );
  OAI22D1BWP U9773 ( .A1(n3680), .A2(n5616), .B1(n4670), .B2(op1[9]), .ZN(
        n6071) );
  AOI22D1BWP U9774 ( .A1(op1[9]), .A2(n4833), .B1(n4654), .B2(n3680), .ZN(
        \mult_x_153/n117 ) );
  AOI22D1BWP U9775 ( .A1(op1[9]), .A2(n5569), .B1(n4667), .B2(n3680), .ZN(
        \mult_x_153/n119 ) );
  AOI22D1BWP U9776 ( .A1(op1[3]), .A2(op2[6]), .B1(n4663), .B2(n5561), .ZN(
        n4824) );
  AOI21D1BWP U9777 ( .A1(n4768), .A2(n5566), .B(n5572), .ZN(n5557) );
  OAI22D1BWP U9778 ( .A1(n6070), .A2(op1[2]), .B1(n4669), .B2(op1[1]), .ZN(
        n5572) );
  AOI22D1BWP U9779 ( .A1(op1[3]), .A2(n5615), .B1(op2[5]), .B2(n5561), .ZN(
        n4825) );
  AOI22D1BWP U9780 ( .A1(op1[7]), .A2(op2[3]), .B1(n5569), .B2(n5605), .ZN(
        n4805) );
  OAI22D1BWP U9781 ( .A1(n4808), .A2(n4802), .B1(n4803), .B2(n4804), .ZN(
        \mult_x_153/n142 ) );
  AOI22D1BWP U9782 ( .A1(op1[7]), .A2(n4663), .B1(op2[6]), .B2(n5605), .ZN(
        n4802) );
  OAI22D1BWP U9783 ( .A1(n4820), .A2(n4813), .B1(n4816), .B2(n4853), .ZN(
        \mult_x_153/n155 ) );
  OAI22D1BWP U9784 ( .A1(n4832), .A2(n5615), .B1(op2[5]), .B2(op1[5]), .ZN(
        n4853) );
  OAI32D1BWP U9785 ( .A1(n4815), .A2(op1[4]), .A3(n4832), .B1(n4809), .B2(
        n4815), .ZN(n4817) );
  AOI22D1BWP U9786 ( .A1(op1[5]), .A2(n4663), .B1(op2[6]), .B2(n4832), .ZN(
        n4813) );
  AOI22D1BWP U9787 ( .A1(op1[9]), .A2(op2[6]), .B1(n4663), .B2(n3680), .ZN(
        n4790) );
  AOI22D1BWP U9788 ( .A1(op1[9]), .A2(n5615), .B1(op2[5]), .B2(n3680), .ZN(
        n4791) );
  OAI22D1BWP U9789 ( .A1(n4808), .A2(n4804), .B1(n4803), .B2(n4807), .ZN(
        \mult_x_153/n143 ) );
  AOI22D1BWP U9790 ( .A1(op1[7]), .A2(n4667), .B1(op2[4]), .B2(n5605), .ZN(
        n4807) );
  OAI32D1BWP U9791 ( .A1(n4800), .A2(op1[6]), .A3(n5605), .B1(n4798), .B2(
        n4800), .ZN(n4806) );
  AOI22D1BWP U9792 ( .A1(op1[7]), .A2(n5615), .B1(op2[5]), .B2(n5605), .ZN(
        n4804) );
  AOI22D1BWP U9793 ( .A1(n4800), .A2(n5605), .B1(n4798), .B2(n4808), .ZN(
        \mult_x_153/n137 ) );
  AOI21D1BWP U9794 ( .A1(n4776), .A2(n4775), .B(\mult_x_153/n88 ), .ZN(
        \mult_x_153/n89 ) );
  NR2XD0BWP U9795 ( .A1(n4775), .A2(n4776), .ZN(\mult_x_153/n88 ) );
  ND3D1BWP U9796 ( .A1(op1[9]), .A2(n5604), .A3(n4782), .ZN(n4775) );
  AOI221D1BWP U9797 ( .A1(n4653), .A2(n3680), .B1(op1[8]), .B2(op1[9]), .C(
        n5555), .ZN(n4796) );
  AOI21D1BWP U9798 ( .A1(op1[9]), .A2(n4680), .B(\mult_x_153/n122 ), .ZN(n4774) );
  NR2XD0BWP U9799 ( .A1(n4680), .A2(op1[9]), .ZN(\mult_x_153/n122 ) );
  AOI22D1BWP U9800 ( .A1(op1[9]), .A2(op2[1]), .B1(n5616), .B2(n3680), .ZN(
        n4795) );
  ND2D1BWP U9801 ( .A1(op1[8]), .A2(op1[7]), .ZN(n5604) );
  OAI21D1BWP U9802 ( .A1(op2[5]), .A2(n5564), .B(n4831), .ZN(\mult_x_153/n181 ) );
  AOI22D1BWP U9803 ( .A1(op2[6]), .A2(n5570), .B1(\mult_x_153/n176 ), .B2(
        n4663), .ZN(n4831) );
  AO222D1BWP U9804 ( .A1(vectorData2[6]), .A2(n4570), .B1(WR), .B2(n5951), 
        .C1(scalarData2[6]), .C2(n4569), .Z(dataOut[6]) );
  ND4D1BWP U9805 ( .A1(n8238), .A2(n8239), .A3(n8240), .A4(n8241), .ZN(
        scalarData2[6]) );
  AOI22D1BWP U9806 ( .A1(n8212), .A2(\srf/regTable[5][6] ), .B1(n8213), .B2(
        \srf/regTable[7][6] ), .ZN(n8241) );
  AOI22D1BWP U9807 ( .A1(n8210), .A2(\srf/regTable[4][6] ), .B1(n8211), .B2(
        \srf/regTable[6][6] ), .ZN(n8240) );
  AOI22D1BWP U9808 ( .A1(n8207), .A2(\srf/regTable[1][6] ), .B1(n8209), .B2(
        \srf/regTable[3][6] ), .ZN(n8239) );
  AOI22D1BWP U9809 ( .A1(n8203), .A2(\srf/regTable[0][6] ), .B1(n8205), .B2(
        \srf/regTable[2][6] ), .ZN(n8238) );
  ND3D1BWP U9810 ( .A1(n5950), .A2(n5949), .A3(n5948), .ZN(n5951) );
  AOI211XD0BWP U9811 ( .A1(n5985), .A2(vectorData2[38]), .B(n5947), .C(n5946), 
        .ZN(n5948) );
  ND4D1BWP U9812 ( .A1(n5945), .A2(n5944), .A3(n5943), .A4(n5942), .ZN(n5946)
         );
  AOI22D1BWP U9813 ( .A1(n5992), .A2(vectorData2[230]), .B1(n5977), .B2(
        vectorData2[134]), .ZN(n5942) );
  ND4D1BWP U9814 ( .A1(n6620), .A2(n6621), .A3(n6622), .A4(n6623), .ZN(
        vectorData2[134]) );
  AOI22D1BWP U9815 ( .A1(n3569), .A2(\vrf/regTable[5][134] ), .B1(n3592), .B2(
        \vrf/regTable[7][134] ), .ZN(n6623) );
  AOI22D1BWP U9816 ( .A1(n3577), .A2(\vrf/regTable[4][134] ), .B1(n3591), .B2(
        \vrf/regTable[6][134] ), .ZN(n6622) );
  AOI22D1BWP U9817 ( .A1(n3571), .A2(\vrf/regTable[1][134] ), .B1(n3568), .B2(
        \vrf/regTable[3][134] ), .ZN(n6621) );
  AOI22D1BWP U9818 ( .A1(n3580), .A2(\vrf/regTable[0][134] ), .B1(n3566), .B2(
        \vrf/regTable[2][134] ), .ZN(n6620) );
  ND4D1BWP U9819 ( .A1(n7004), .A2(n7005), .A3(n7006), .A4(n7007), .ZN(
        vectorData2[230]) );
  AOI22D1BWP U9820 ( .A1(n3569), .A2(\vrf/regTable[5][230] ), .B1(n3592), .B2(
        \vrf/regTable[7][230] ), .ZN(n7007) );
  AOI22D1BWP U9821 ( .A1(n3577), .A2(\vrf/regTable[4][230] ), .B1(n3591), .B2(
        \vrf/regTable[6][230] ), .ZN(n7006) );
  AOI22D1BWP U9822 ( .A1(n3571), .A2(\vrf/regTable[1][230] ), .B1(n3568), .B2(
        \vrf/regTable[3][230] ), .ZN(n7005) );
  AOI22D1BWP U9823 ( .A1(n3580), .A2(\vrf/regTable[0][230] ), .B1(n3566), .B2(
        \vrf/regTable[2][230] ), .ZN(n7004) );
  AOI22D1BWP U9824 ( .A1(n5974), .A2(vectorData2[54]), .B1(n5972), .B2(
        vectorData2[118]), .ZN(n5943) );
  ND4D1BWP U9825 ( .A1(n6556), .A2(n6557), .A3(n6558), .A4(n6559), .ZN(
        vectorData2[118]) );
  AOI22D1BWP U9826 ( .A1(n3569), .A2(\vrf/regTable[5][118] ), .B1(n3578), .B2(
        \vrf/regTable[7][118] ), .ZN(n6559) );
  AOI22D1BWP U9827 ( .A1(n3577), .A2(\vrf/regTable[4][118] ), .B1(n3573), .B2(
        \vrf/regTable[6][118] ), .ZN(n6558) );
  AOI22D1BWP U9828 ( .A1(n3571), .A2(\vrf/regTable[1][118] ), .B1(n3597), .B2(
        \vrf/regTable[3][118] ), .ZN(n6557) );
  AOI22D1BWP U9829 ( .A1(n3580), .A2(\vrf/regTable[0][118] ), .B1(n3593), .B2(
        \vrf/regTable[2][118] ), .ZN(n6556) );
  ND4D1BWP U9830 ( .A1(n6300), .A2(n6301), .A3(n6302), .A4(n6303), .ZN(
        vectorData2[54]) );
  AOI22D1BWP U9831 ( .A1(n3569), .A2(\vrf/regTable[5][54] ), .B1(n3592), .B2(
        \vrf/regTable[7][54] ), .ZN(n6303) );
  AOI22D1BWP U9832 ( .A1(n3577), .A2(\vrf/regTable[4][54] ), .B1(n3591), .B2(
        \vrf/regTable[6][54] ), .ZN(n6302) );
  AOI22D1BWP U9833 ( .A1(n3571), .A2(\vrf/regTable[1][54] ), .B1(n3568), .B2(
        \vrf/regTable[3][54] ), .ZN(n6301) );
  AOI22D1BWP U9834 ( .A1(n3580), .A2(\vrf/regTable[0][54] ), .B1(n3566), .B2(
        \vrf/regTable[2][54] ), .ZN(n6300) );
  AOI22D1BWP U9835 ( .A1(n5973), .A2(vectorData2[70]), .B1(n5983), .B2(
        vectorData2[150]), .ZN(n5944) );
  ND4D1BWP U9836 ( .A1(n6684), .A2(n6685), .A3(n6686), .A4(n6687), .ZN(
        vectorData2[150]) );
  AOI22D1BWP U9837 ( .A1(n3569), .A2(\vrf/regTable[5][150] ), .B1(n3578), .B2(
        \vrf/regTable[7][150] ), .ZN(n6687) );
  AOI22D1BWP U9838 ( .A1(n3577), .A2(\vrf/regTable[4][150] ), .B1(n3573), .B2(
        \vrf/regTable[6][150] ), .ZN(n6686) );
  AOI22D1BWP U9839 ( .A1(n3571), .A2(\vrf/regTable[1][150] ), .B1(n3597), .B2(
        \vrf/regTable[3][150] ), .ZN(n6685) );
  AOI22D1BWP U9840 ( .A1(n3580), .A2(\vrf/regTable[0][150] ), .B1(n3593), .B2(
        \vrf/regTable[2][150] ), .ZN(n6684) );
  ND4D1BWP U9841 ( .A1(n6364), .A2(n6365), .A3(n6366), .A4(n6367), .ZN(
        vectorData2[70]) );
  AOI22D1BWP U9842 ( .A1(n3569), .A2(\vrf/regTable[5][70] ), .B1(n3578), .B2(
        \vrf/regTable[7][70] ), .ZN(n6367) );
  AOI22D1BWP U9843 ( .A1(n3577), .A2(\vrf/regTable[4][70] ), .B1(n3573), .B2(
        \vrf/regTable[6][70] ), .ZN(n6366) );
  AOI22D1BWP U9844 ( .A1(n3571), .A2(\vrf/regTable[1][70] ), .B1(n3597), .B2(
        \vrf/regTable[3][70] ), .ZN(n6365) );
  AOI22D1BWP U9845 ( .A1(n3580), .A2(\vrf/regTable[0][70] ), .B1(n3593), .B2(
        \vrf/regTable[2][70] ), .ZN(n6364) );
  AOI22D1BWP U9846 ( .A1(n5978), .A2(vectorData2[198]), .B1(n5982), .B2(
        vectorData2[22]), .ZN(n5945) );
  ND4D1BWP U9847 ( .A1(n6172), .A2(n6173), .A3(n6174), .A4(n6175), .ZN(
        vectorData2[22]) );
  AOI22D1BWP U9848 ( .A1(n6082), .A2(\vrf/regTable[5][22] ), .B1(n3592), .B2(
        \vrf/regTable[7][22] ), .ZN(n6175) );
  AOI22D1BWP U9849 ( .A1(n3577), .A2(\vrf/regTable[4][22] ), .B1(n3591), .B2(
        \vrf/regTable[6][22] ), .ZN(n6174) );
  AOI22D1BWP U9850 ( .A1(n6077), .A2(\vrf/regTable[1][22] ), .B1(n3568), .B2(
        \vrf/regTable[3][22] ), .ZN(n6173) );
  AOI22D1BWP U9851 ( .A1(n3580), .A2(\vrf/regTable[0][22] ), .B1(n3566), .B2(
        \vrf/regTable[2][22] ), .ZN(n6172) );
  ND4D1BWP U9852 ( .A1(n6876), .A2(n6877), .A3(n6878), .A4(n6879), .ZN(
        vectorData2[198]) );
  AOI22D1BWP U9853 ( .A1(n3569), .A2(\vrf/regTable[5][198] ), .B1(n3578), .B2(
        \vrf/regTable[7][198] ), .ZN(n6879) );
  AOI22D1BWP U9854 ( .A1(n3577), .A2(\vrf/regTable[4][198] ), .B1(n3573), .B2(
        \vrf/regTable[6][198] ), .ZN(n6878) );
  AOI22D1BWP U9855 ( .A1(n3571), .A2(\vrf/regTable[1][198] ), .B1(n3597), .B2(
        \vrf/regTable[3][198] ), .ZN(n6877) );
  AOI22D1BWP U9856 ( .A1(n3580), .A2(\vrf/regTable[0][198] ), .B1(n3593), .B2(
        \vrf/regTable[2][198] ), .ZN(n6876) );
  AO22D1BWP U9857 ( .A1(n5979), .A2(vectorData2[86]), .B1(n5976), .B2(
        vectorData2[102]), .Z(n5947) );
  ND4D1BWP U9858 ( .A1(n6492), .A2(n6493), .A3(n6494), .A4(n6495), .ZN(
        vectorData2[102]) );
  AOI22D1BWP U9859 ( .A1(n3569), .A2(\vrf/regTable[5][102] ), .B1(n3578), .B2(
        \vrf/regTable[7][102] ), .ZN(n6495) );
  AOI22D1BWP U9860 ( .A1(n3577), .A2(\vrf/regTable[4][102] ), .B1(n3573), .B2(
        \vrf/regTable[6][102] ), .ZN(n6494) );
  AOI22D1BWP U9861 ( .A1(n3571), .A2(\vrf/regTable[1][102] ), .B1(n3597), .B2(
        \vrf/regTable[3][102] ), .ZN(n6493) );
  AOI22D1BWP U9862 ( .A1(n3580), .A2(\vrf/regTable[0][102] ), .B1(n3593), .B2(
        \vrf/regTable[2][102] ), .ZN(n6492) );
  ND4D1BWP U9863 ( .A1(n6428), .A2(n6429), .A3(n6430), .A4(n6431), .ZN(
        vectorData2[86]) );
  AOI22D1BWP U9864 ( .A1(n3569), .A2(\vrf/regTable[5][86] ), .B1(n3592), .B2(
        \vrf/regTable[7][86] ), .ZN(n6431) );
  AOI22D1BWP U9865 ( .A1(n8210), .A2(\vrf/regTable[4][86] ), .B1(n3591), .B2(
        \vrf/regTable[6][86] ), .ZN(n6430) );
  AOI22D1BWP U9866 ( .A1(n3571), .A2(\vrf/regTable[1][86] ), .B1(n3568), .B2(
        \vrf/regTable[3][86] ), .ZN(n6429) );
  AOI22D1BWP U9867 ( .A1(n8203), .A2(\vrf/regTable[0][86] ), .B1(n3566), .B2(
        \vrf/regTable[2][86] ), .ZN(n6428) );
  ND4D1BWP U9868 ( .A1(n6236), .A2(n6237), .A3(n6238), .A4(n6239), .ZN(
        vectorData2[38]) );
  AOI22D1BWP U9869 ( .A1(n6082), .A2(\vrf/regTable[5][38] ), .B1(n3578), .B2(
        \vrf/regTable[7][38] ), .ZN(n6239) );
  AOI22D1BWP U9870 ( .A1(n3577), .A2(\vrf/regTable[4][38] ), .B1(n3573), .B2(
        \vrf/regTable[6][38] ), .ZN(n6238) );
  AOI22D1BWP U9871 ( .A1(n6077), .A2(\vrf/regTable[1][38] ), .B1(n3597), .B2(
        \vrf/regTable[3][38] ), .ZN(n6237) );
  AOI22D1BWP U9872 ( .A1(n3580), .A2(\vrf/regTable[0][38] ), .B1(n3593), .B2(
        \vrf/regTable[2][38] ), .ZN(n6236) );
  AOI22D1BWP U9873 ( .A1(n5981), .A2(vectorData2[182]), .B1(n5975), .B2(
        vectorData2[166]), .ZN(n5949) );
  ND4D1BWP U9874 ( .A1(n6748), .A2(n6749), .A3(n6750), .A4(n6751), .ZN(
        vectorData2[166]) );
  AOI22D1BWP U9875 ( .A1(n3569), .A2(\vrf/regTable[5][166] ), .B1(n3592), .B2(
        \vrf/regTable[7][166] ), .ZN(n6751) );
  AOI22D1BWP U9876 ( .A1(n3577), .A2(\vrf/regTable[4][166] ), .B1(n3591), .B2(
        \vrf/regTable[6][166] ), .ZN(n6750) );
  AOI22D1BWP U9877 ( .A1(n3571), .A2(\vrf/regTable[1][166] ), .B1(n3568), .B2(
        \vrf/regTable[3][166] ), .ZN(n6749) );
  AOI22D1BWP U9878 ( .A1(n3580), .A2(\vrf/regTable[0][166] ), .B1(n3566), .B2(
        \vrf/regTable[2][166] ), .ZN(n6748) );
  ND4D1BWP U9879 ( .A1(n6812), .A2(n6813), .A3(n6814), .A4(n6815), .ZN(
        vectorData2[182]) );
  AOI22D1BWP U9880 ( .A1(n3569), .A2(\vrf/regTable[5][182] ), .B1(n3592), .B2(
        \vrf/regTable[7][182] ), .ZN(n6815) );
  AOI22D1BWP U9881 ( .A1(n3577), .A2(\vrf/regTable[4][182] ), .B1(n3591), .B2(
        \vrf/regTable[6][182] ), .ZN(n6814) );
  AOI22D1BWP U9882 ( .A1(n3571), .A2(\vrf/regTable[1][182] ), .B1(n3568), .B2(
        \vrf/regTable[3][182] ), .ZN(n6813) );
  AOI22D1BWP U9883 ( .A1(n3580), .A2(\vrf/regTable[0][182] ), .B1(n3566), .B2(
        \vrf/regTable[2][182] ), .ZN(n6812) );
  AOI22D1BWP U9884 ( .A1(n5984), .A2(vectorData2[214]), .B1(n5980), .B2(
        vectorData2[246]), .ZN(n5950) );
  ND4D1BWP U9885 ( .A1(n7068), .A2(n7069), .A3(n7070), .A4(n7071), .ZN(
        vectorData2[246]) );
  AOI22D1BWP U9886 ( .A1(n6082), .A2(\vrf/regTable[5][246] ), .B1(n3578), .B2(
        \vrf/regTable[7][246] ), .ZN(n7071) );
  AOI22D1BWP U9887 ( .A1(n3577), .A2(\vrf/regTable[4][246] ), .B1(n3573), .B2(
        \vrf/regTable[6][246] ), .ZN(n7070) );
  AOI22D1BWP U9888 ( .A1(n6077), .A2(\vrf/regTable[1][246] ), .B1(n3597), .B2(
        \vrf/regTable[3][246] ), .ZN(n7069) );
  AOI22D1BWP U9889 ( .A1(n3580), .A2(\vrf/regTable[0][246] ), .B1(n3593), .B2(
        \vrf/regTable[2][246] ), .ZN(n7068) );
  ND4D1BWP U9890 ( .A1(n6940), .A2(n6941), .A3(n6942), .A4(n6943), .ZN(
        vectorData2[214]) );
  AOI22D1BWP U9891 ( .A1(n6082), .A2(\vrf/regTable[5][214] ), .B1(n3578), .B2(
        \vrf/regTable[7][214] ), .ZN(n6943) );
  AOI22D1BWP U9892 ( .A1(n3577), .A2(\vrf/regTable[4][214] ), .B1(n3573), .B2(
        \vrf/regTable[6][214] ), .ZN(n6942) );
  AOI22D1BWP U9893 ( .A1(n6077), .A2(\vrf/regTable[1][214] ), .B1(n3597), .B2(
        \vrf/regTable[3][214] ), .ZN(n6941) );
  AOI22D1BWP U9894 ( .A1(n3580), .A2(\vrf/regTable[0][214] ), .B1(n3593), .B2(
        \vrf/regTable[2][214] ), .ZN(n6940) );
  ND4D1BWP U9895 ( .A1(n6108), .A2(n6109), .A3(n6110), .A4(n6111), .ZN(
        vectorData2[6]) );
  AOI22D1BWP U9896 ( .A1(n3569), .A2(\vrf/regTable[5][6] ), .B1(n3592), .B2(
        \vrf/regTable[7][6] ), .ZN(n6111) );
  AOI22D1BWP U9897 ( .A1(n3577), .A2(\vrf/regTable[4][6] ), .B1(n3591), .B2(
        \vrf/regTable[6][6] ), .ZN(n6110) );
  AOI22D1BWP U9898 ( .A1(n3571), .A2(\vrf/regTable[1][6] ), .B1(n3568), .B2(
        \vrf/regTable[3][6] ), .ZN(n6109) );
  AOI22D1BWP U9899 ( .A1(n3580), .A2(\vrf/regTable[0][6] ), .B1(n3566), .B2(
        \vrf/regTable[2][6] ), .ZN(n6108) );
  AO222D1BWP U9900 ( .A1(WR), .A2(n5931), .B1(n4570), .B2(vectorData2[4]), 
        .C1(n4569), .C2(scalarData2[4]), .Z(dataOut[4]) );
  ND4D1BWP U9901 ( .A1(n8230), .A2(n8231), .A3(n8232), .A4(n8233), .ZN(
        scalarData2[4]) );
  AOI22D1BWP U9902 ( .A1(n8212), .A2(\srf/regTable[5][4] ), .B1(n8213), .B2(
        \srf/regTable[7][4] ), .ZN(n8233) );
  AOI22D1BWP U9903 ( .A1(n8210), .A2(\srf/regTable[4][4] ), .B1(n8211), .B2(
        \srf/regTable[6][4] ), .ZN(n8232) );
  AOI22D1BWP U9904 ( .A1(n8207), .A2(\srf/regTable[1][4] ), .B1(n8209), .B2(
        \srf/regTable[3][4] ), .ZN(n8231) );
  AOI22D1BWP U9905 ( .A1(n8203), .A2(\srf/regTable[0][4] ), .B1(n8205), .B2(
        \srf/regTable[2][4] ), .ZN(n8230) );
  ND4D1BWP U9906 ( .A1(n6100), .A2(n6101), .A3(n6102), .A4(n6103), .ZN(
        vectorData2[4]) );
  AOI22D1BWP U9907 ( .A1(n3569), .A2(\vrf/regTable[5][4] ), .B1(n3578), .B2(
        \vrf/regTable[7][4] ), .ZN(n6103) );
  AOI22D1BWP U9908 ( .A1(n3577), .A2(\vrf/regTable[4][4] ), .B1(n3573), .B2(
        \vrf/regTable[6][4] ), .ZN(n6102) );
  AOI22D1BWP U9909 ( .A1(n3571), .A2(\vrf/regTable[1][4] ), .B1(n3597), .B2(
        \vrf/regTable[3][4] ), .ZN(n6101) );
  AOI22D1BWP U9910 ( .A1(n3580), .A2(\vrf/regTable[0][4] ), .B1(n3593), .B2(
        \vrf/regTable[2][4] ), .ZN(n6100) );
  ND3D1BWP U9911 ( .A1(n5930), .A2(n5929), .A3(n5928), .ZN(n5931) );
  AOI211XD0BWP U9912 ( .A1(n5985), .A2(vectorData2[36]), .B(n5927), .C(n5926), 
        .ZN(n5928) );
  ND4D1BWP U9913 ( .A1(n5925), .A2(n5924), .A3(n5923), .A4(n5922), .ZN(n5926)
         );
  AOI22D1BWP U9914 ( .A1(n5982), .A2(vectorData2[20]), .B1(n5976), .B2(
        vectorData2[100]), .ZN(n5922) );
  ND4D1BWP U9915 ( .A1(n6484), .A2(n6485), .A3(n6486), .A4(n6487), .ZN(
        vectorData2[100]) );
  AOI22D1BWP U9916 ( .A1(n3569), .A2(\vrf/regTable[5][100] ), .B1(n3578), .B2(
        \vrf/regTable[7][100] ), .ZN(n6487) );
  AOI22D1BWP U9917 ( .A1(n3577), .A2(\vrf/regTable[4][100] ), .B1(n3573), .B2(
        \vrf/regTable[6][100] ), .ZN(n6486) );
  AOI22D1BWP U9918 ( .A1(n3571), .A2(\vrf/regTable[1][100] ), .B1(n3597), .B2(
        \vrf/regTable[3][100] ), .ZN(n6485) );
  AOI22D1BWP U9919 ( .A1(n3580), .A2(\vrf/regTable[0][100] ), .B1(n3593), .B2(
        \vrf/regTable[2][100] ), .ZN(n6484) );
  ND4D1BWP U9920 ( .A1(n6164), .A2(n6165), .A3(n6166), .A4(n6167), .ZN(
        vectorData2[20]) );
  AOI22D1BWP U9921 ( .A1(n3569), .A2(\vrf/regTable[5][20] ), .B1(n3592), .B2(
        \vrf/regTable[7][20] ), .ZN(n6167) );
  AOI22D1BWP U9922 ( .A1(n3577), .A2(\vrf/regTable[4][20] ), .B1(n3591), .B2(
        \vrf/regTable[6][20] ), .ZN(n6166) );
  AOI22D1BWP U9923 ( .A1(n3571), .A2(\vrf/regTable[1][20] ), .B1(n3568), .B2(
        \vrf/regTable[3][20] ), .ZN(n6165) );
  AOI22D1BWP U9924 ( .A1(n3580), .A2(\vrf/regTable[0][20] ), .B1(n3566), .B2(
        \vrf/regTable[2][20] ), .ZN(n6164) );
  AOI22D1BWP U9925 ( .A1(n5981), .A2(vectorData2[180]), .B1(n5974), .B2(
        vectorData2[52]), .ZN(n5923) );
  ND4D1BWP U9926 ( .A1(n6292), .A2(n6293), .A3(n6294), .A4(n6295), .ZN(
        vectorData2[52]) );
  AOI22D1BWP U9927 ( .A1(n3569), .A2(\vrf/regTable[5][52] ), .B1(n3592), .B2(
        \vrf/regTable[7][52] ), .ZN(n6295) );
  AOI22D1BWP U9928 ( .A1(n3577), .A2(\vrf/regTable[4][52] ), .B1(n3591), .B2(
        \vrf/regTable[6][52] ), .ZN(n6294) );
  AOI22D1BWP U9929 ( .A1(n3571), .A2(\vrf/regTable[1][52] ), .B1(n3568), .B2(
        \vrf/regTable[3][52] ), .ZN(n6293) );
  AOI22D1BWP U9930 ( .A1(n3580), .A2(\vrf/regTable[0][52] ), .B1(n3566), .B2(
        \vrf/regTable[2][52] ), .ZN(n6292) );
  ND4D1BWP U9931 ( .A1(n6804), .A2(n6805), .A3(n6806), .A4(n6807), .ZN(
        vectorData2[180]) );
  AOI22D1BWP U9932 ( .A1(n3569), .A2(\vrf/regTable[5][180] ), .B1(n3592), .B2(
        \vrf/regTable[7][180] ), .ZN(n6807) );
  AOI22D1BWP U9933 ( .A1(n3577), .A2(\vrf/regTable[4][180] ), .B1(n3591), .B2(
        \vrf/regTable[6][180] ), .ZN(n6806) );
  AOI22D1BWP U9934 ( .A1(n3571), .A2(\vrf/regTable[1][180] ), .B1(n3568), .B2(
        \vrf/regTable[3][180] ), .ZN(n6805) );
  AOI22D1BWP U9935 ( .A1(n3580), .A2(\vrf/regTable[0][180] ), .B1(n3566), .B2(
        \vrf/regTable[2][180] ), .ZN(n6804) );
  AOI22D1BWP U9936 ( .A1(n5978), .A2(vectorData2[196]), .B1(n5973), .B2(
        vectorData2[68]), .ZN(n5924) );
  ND4D1BWP U9937 ( .A1(n6356), .A2(n6357), .A3(n6358), .A4(n6359), .ZN(
        vectorData2[68]) );
  AOI22D1BWP U9938 ( .A1(n3569), .A2(\vrf/regTable[5][68] ), .B1(n3592), .B2(
        \vrf/regTable[7][68] ), .ZN(n6359) );
  AOI22D1BWP U9939 ( .A1(n3577), .A2(\vrf/regTable[4][68] ), .B1(n3591), .B2(
        \vrf/regTable[6][68] ), .ZN(n6358) );
  AOI22D1BWP U9940 ( .A1(n3571), .A2(\vrf/regTable[1][68] ), .B1(n3568), .B2(
        \vrf/regTable[3][68] ), .ZN(n6357) );
  AOI22D1BWP U9941 ( .A1(n3580), .A2(\vrf/regTable[0][68] ), .B1(n3566), .B2(
        \vrf/regTable[2][68] ), .ZN(n6356) );
  ND4D1BWP U9942 ( .A1(n6868), .A2(n6869), .A3(n6870), .A4(n6871), .ZN(
        vectorData2[196]) );
  AOI22D1BWP U9943 ( .A1(n3569), .A2(\vrf/regTable[5][196] ), .B1(n3578), .B2(
        \vrf/regTable[7][196] ), .ZN(n6871) );
  AOI22D1BWP U9944 ( .A1(n3577), .A2(\vrf/regTable[4][196] ), .B1(n3573), .B2(
        \vrf/regTable[6][196] ), .ZN(n6870) );
  AOI22D1BWP U9945 ( .A1(n3571), .A2(\vrf/regTable[1][196] ), .B1(n3597), .B2(
        \vrf/regTable[3][196] ), .ZN(n6869) );
  AOI22D1BWP U9946 ( .A1(n3580), .A2(\vrf/regTable[0][196] ), .B1(n3593), .B2(
        \vrf/regTable[2][196] ), .ZN(n6868) );
  AOI22D1BWP U9947 ( .A1(n5992), .A2(vectorData2[228]), .B1(n5975), .B2(
        vectorData2[164]), .ZN(n5925) );
  ND4D1BWP U9948 ( .A1(n6740), .A2(n6741), .A3(n6742), .A4(n6743), .ZN(
        vectorData2[164]) );
  AOI22D1BWP U9949 ( .A1(n3569), .A2(\vrf/regTable[5][164] ), .B1(n3578), .B2(
        \vrf/regTable[7][164] ), .ZN(n6743) );
  AOI22D1BWP U9950 ( .A1(n3577), .A2(\vrf/regTable[4][164] ), .B1(n3573), .B2(
        \vrf/regTable[6][164] ), .ZN(n6742) );
  AOI22D1BWP U9951 ( .A1(n3571), .A2(\vrf/regTable[1][164] ), .B1(n3597), .B2(
        \vrf/regTable[3][164] ), .ZN(n6741) );
  AOI22D1BWP U9952 ( .A1(n3580), .A2(\vrf/regTable[0][164] ), .B1(n3593), .B2(
        \vrf/regTable[2][164] ), .ZN(n6740) );
  ND4D1BWP U9953 ( .A1(n6996), .A2(n6997), .A3(n6998), .A4(n6999), .ZN(
        vectorData2[228]) );
  AOI22D1BWP U9954 ( .A1(n3569), .A2(\vrf/regTable[5][228] ), .B1(n3578), .B2(
        \vrf/regTable[7][228] ), .ZN(n6999) );
  AOI22D1BWP U9955 ( .A1(n3577), .A2(\vrf/regTable[4][228] ), .B1(n3573), .B2(
        \vrf/regTable[6][228] ), .ZN(n6998) );
  AOI22D1BWP U9956 ( .A1(n3571), .A2(\vrf/regTable[1][228] ), .B1(n3597), .B2(
        \vrf/regTable[3][228] ), .ZN(n6997) );
  AOI22D1BWP U9957 ( .A1(n3580), .A2(\vrf/regTable[0][228] ), .B1(n3593), .B2(
        \vrf/regTable[2][228] ), .ZN(n6996) );
  AO22D1BWP U9958 ( .A1(n5979), .A2(vectorData2[84]), .B1(n5977), .B2(
        vectorData2[132]), .Z(n5927) );
  ND4D1BWP U9959 ( .A1(n6612), .A2(n6613), .A3(n6614), .A4(n6615), .ZN(
        vectorData2[132]) );
  AOI22D1BWP U9960 ( .A1(n3569), .A2(\vrf/regTable[5][132] ), .B1(n3592), .B2(
        \vrf/regTable[7][132] ), .ZN(n6615) );
  AOI22D1BWP U9961 ( .A1(n3577), .A2(\vrf/regTable[4][132] ), .B1(n3591), .B2(
        \vrf/regTable[6][132] ), .ZN(n6614) );
  AOI22D1BWP U9962 ( .A1(n3571), .A2(\vrf/regTable[1][132] ), .B1(n3568), .B2(
        \vrf/regTable[3][132] ), .ZN(n6613) );
  AOI22D1BWP U9963 ( .A1(n3580), .A2(\vrf/regTable[0][132] ), .B1(n3566), .B2(
        \vrf/regTable[2][132] ), .ZN(n6612) );
  ND4D1BWP U9964 ( .A1(n6420), .A2(n6421), .A3(n6422), .A4(n6423), .ZN(
        vectorData2[84]) );
  AOI22D1BWP U9965 ( .A1(n6082), .A2(\vrf/regTable[5][84] ), .B1(n3592), .B2(
        \vrf/regTable[7][84] ), .ZN(n6423) );
  AOI22D1BWP U9966 ( .A1(n3577), .A2(\vrf/regTable[4][84] ), .B1(n3591), .B2(
        \vrf/regTable[6][84] ), .ZN(n6422) );
  AOI22D1BWP U9967 ( .A1(n6077), .A2(\vrf/regTable[1][84] ), .B1(n3568), .B2(
        \vrf/regTable[3][84] ), .ZN(n6421) );
  AOI22D1BWP U9968 ( .A1(n3580), .A2(\vrf/regTable[0][84] ), .B1(n3566), .B2(
        \vrf/regTable[2][84] ), .ZN(n6420) );
  ND4D1BWP U9969 ( .A1(n6228), .A2(n6229), .A3(n6230), .A4(n6231), .ZN(
        vectorData2[36]) );
  AOI22D1BWP U9970 ( .A1(n3569), .A2(\vrf/regTable[5][36] ), .B1(n3592), .B2(
        \vrf/regTable[7][36] ), .ZN(n6231) );
  AOI22D1BWP U9971 ( .A1(n8210), .A2(\vrf/regTable[4][36] ), .B1(n3591), .B2(
        \vrf/regTable[6][36] ), .ZN(n6230) );
  AOI22D1BWP U9972 ( .A1(n3571), .A2(\vrf/regTable[1][36] ), .B1(n3568), .B2(
        \vrf/regTable[3][36] ), .ZN(n6229) );
  AOI22D1BWP U9973 ( .A1(n8203), .A2(\vrf/regTable[0][36] ), .B1(n3566), .B2(
        \vrf/regTable[2][36] ), .ZN(n6228) );
  AOI22D1BWP U9974 ( .A1(n5984), .A2(vectorData2[212]), .B1(n5972), .B2(
        vectorData2[116]), .ZN(n5929) );
  ND4D1BWP U9975 ( .A1(n6548), .A2(n6549), .A3(n6550), .A4(n6551), .ZN(
        vectorData2[116]) );
  AOI22D1BWP U9976 ( .A1(n6082), .A2(\vrf/regTable[5][116] ), .B1(n3578), .B2(
        \vrf/regTable[7][116] ), .ZN(n6551) );
  AOI22D1BWP U9977 ( .A1(n3577), .A2(\vrf/regTable[4][116] ), .B1(n3573), .B2(
        \vrf/regTable[6][116] ), .ZN(n6550) );
  AOI22D1BWP U9978 ( .A1(n6077), .A2(\vrf/regTable[1][116] ), .B1(n3597), .B2(
        \vrf/regTable[3][116] ), .ZN(n6549) );
  AOI22D1BWP U9979 ( .A1(n3580), .A2(\vrf/regTable[0][116] ), .B1(n3593), .B2(
        \vrf/regTable[2][116] ), .ZN(n6548) );
  ND4D1BWP U9980 ( .A1(n6932), .A2(n6933), .A3(n6934), .A4(n6935), .ZN(
        vectorData2[212]) );
  AOI22D1BWP U9981 ( .A1(n6082), .A2(\vrf/regTable[5][212] ), .B1(n3592), .B2(
        \vrf/regTable[7][212] ), .ZN(n6935) );
  AOI22D1BWP U9982 ( .A1(n3577), .A2(\vrf/regTable[4][212] ), .B1(n3591), .B2(
        \vrf/regTable[6][212] ), .ZN(n6934) );
  AOI22D1BWP U9983 ( .A1(n6077), .A2(\vrf/regTable[1][212] ), .B1(n3568), .B2(
        \vrf/regTable[3][212] ), .ZN(n6933) );
  AOI22D1BWP U9984 ( .A1(n3580), .A2(\vrf/regTable[0][212] ), .B1(n3566), .B2(
        \vrf/regTable[2][212] ), .ZN(n6932) );
  AOI22D1BWP U9985 ( .A1(n5983), .A2(vectorData2[148]), .B1(n5980), .B2(
        vectorData2[244]), .ZN(n5930) );
  ND4D1BWP U9986 ( .A1(n7060), .A2(n7061), .A3(n7062), .A4(n7063), .ZN(
        vectorData2[244]) );
  AOI22D1BWP U9987 ( .A1(n3569), .A2(\vrf/regTable[5][244] ), .B1(n3578), .B2(
        \vrf/regTable[7][244] ), .ZN(n7063) );
  AOI22D1BWP U9988 ( .A1(n3577), .A2(\vrf/regTable[4][244] ), .B1(n3573), .B2(
        \vrf/regTable[6][244] ), .ZN(n7062) );
  AOI22D1BWP U9989 ( .A1(n3571), .A2(\vrf/regTable[1][244] ), .B1(n3597), .B2(
        \vrf/regTable[3][244] ), .ZN(n7061) );
  AOI22D1BWP U9990 ( .A1(n3580), .A2(\vrf/regTable[0][244] ), .B1(n3593), .B2(
        \vrf/regTable[2][244] ), .ZN(n7060) );
  ND4D1BWP U9991 ( .A1(n6676), .A2(n6677), .A3(n6678), .A4(n6679), .ZN(
        vectorData2[148]) );
  AOI22D1BWP U9992 ( .A1(n6082), .A2(\vrf/regTable[5][148] ), .B1(n3578), .B2(
        \vrf/regTable[7][148] ), .ZN(n6679) );
  AOI22D1BWP U9993 ( .A1(n3577), .A2(\vrf/regTable[4][148] ), .B1(n3573), .B2(
        \vrf/regTable[6][148] ), .ZN(n6678) );
  AOI22D1BWP U9994 ( .A1(n6077), .A2(\vrf/regTable[1][148] ), .B1(n3597), .B2(
        \vrf/regTable[3][148] ), .ZN(n6677) );
  AOI22D1BWP U9995 ( .A1(n3580), .A2(\vrf/regTable[0][148] ), .B1(n3593), .B2(
        \vrf/regTable[2][148] ), .ZN(n6676) );
  AO222D1BWP U9996 ( .A1(vectorData2[5]), .A2(n4570), .B1(WR), .B2(n5941), 
        .C1(scalarData2[5]), .C2(n4569), .Z(dataOut[5]) );
  ND4D1BWP U9997 ( .A1(n8234), .A2(n8235), .A3(n8236), .A4(n8237), .ZN(
        scalarData2[5]) );
  AOI22D1BWP U9998 ( .A1(n8212), .A2(\srf/regTable[5][5] ), .B1(n8213), .B2(
        \srf/regTable[7][5] ), .ZN(n8237) );
  AOI22D1BWP U9999 ( .A1(n8210), .A2(\srf/regTable[4][5] ), .B1(n8211), .B2(
        \srf/regTable[6][5] ), .ZN(n8236) );
  AOI22D1BWP U10000 ( .A1(n8207), .A2(\srf/regTable[1][5] ), .B1(n8209), .B2(
        \srf/regTable[3][5] ), .ZN(n8235) );
  AOI22D1BWP U10001 ( .A1(n8203), .A2(\srf/regTable[0][5] ), .B1(n8205), .B2(
        \srf/regTable[2][5] ), .ZN(n8234) );
  ND3D1BWP U10002 ( .A1(n5940), .A2(n5939), .A3(n5938), .ZN(n5941) );
  AOI211XD0BWP U10003 ( .A1(n5979), .A2(vectorData2[85]), .B(n5937), .C(n5936), 
        .ZN(n5938) );
  ND4D1BWP U10004 ( .A1(n5935), .A2(n5934), .A3(n5933), .A4(n5932), .ZN(n5936)
         );
  AOI22D1BWP U10005 ( .A1(n5992), .A2(vectorData2[229]), .B1(n5978), .B2(
        vectorData2[197]), .ZN(n5932) );
  ND4D1BWP U10006 ( .A1(n6872), .A2(n6873), .A3(n6874), .A4(n6875), .ZN(
        vectorData2[197]) );
  AOI22D1BWP U10007 ( .A1(n3569), .A2(\vrf/regTable[5][197] ), .B1(n6083), 
        .B2(\vrf/regTable[7][197] ), .ZN(n6875) );
  AOI22D1BWP U10008 ( .A1(n3577), .A2(\vrf/regTable[4][197] ), .B1(n6081), 
        .B2(\vrf/regTable[6][197] ), .ZN(n6874) );
  AOI22D1BWP U10009 ( .A1(n3571), .A2(\vrf/regTable[1][197] ), .B1(n6079), 
        .B2(\vrf/regTable[3][197] ), .ZN(n6873) );
  AOI22D1BWP U10010 ( .A1(n3580), .A2(\vrf/regTable[0][197] ), .B1(n6075), 
        .B2(\vrf/regTable[2][197] ), .ZN(n6872) );
  ND4D1BWP U10011 ( .A1(n7000), .A2(n7001), .A3(n7002), .A4(n7003), .ZN(
        vectorData2[229]) );
  AOI22D1BWP U10012 ( .A1(n3569), .A2(\vrf/regTable[5][229] ), .B1(n3592), 
        .B2(\vrf/regTable[7][229] ), .ZN(n7003) );
  AOI22D1BWP U10013 ( .A1(n6080), .A2(\vrf/regTable[4][229] ), .B1(n3591), 
        .B2(\vrf/regTable[6][229] ), .ZN(n7002) );
  AOI22D1BWP U10014 ( .A1(n3571), .A2(\vrf/regTable[1][229] ), .B1(n3568), 
        .B2(\vrf/regTable[3][229] ), .ZN(n7001) );
  AOI22D1BWP U10015 ( .A1(n6073), .A2(\vrf/regTable[0][229] ), .B1(n3566), 
        .B2(\vrf/regTable[2][229] ), .ZN(n7000) );
  AOI22D1BWP U10016 ( .A1(n5972), .A2(vectorData2[117]), .B1(n5982), .B2(
        vectorData2[21]), .ZN(n5933) );
  ND4D1BWP U10017 ( .A1(n6168), .A2(n6169), .A3(n6170), .A4(n6171), .ZN(
        vectorData2[21]) );
  AOI22D1BWP U10018 ( .A1(n3569), .A2(\vrf/regTable[5][21] ), .B1(n3578), .B2(
        \vrf/regTable[7][21] ), .ZN(n6171) );
  AOI22D1BWP U10019 ( .A1(n3577), .A2(\vrf/regTable[4][21] ), .B1(n3573), .B2(
        \vrf/regTable[6][21] ), .ZN(n6170) );
  AOI22D1BWP U10020 ( .A1(n3571), .A2(\vrf/regTable[1][21] ), .B1(n3597), .B2(
        \vrf/regTable[3][21] ), .ZN(n6169) );
  AOI22D1BWP U10021 ( .A1(n3580), .A2(\vrf/regTable[0][21] ), .B1(n3593), .B2(
        \vrf/regTable[2][21] ), .ZN(n6168) );
  ND4D1BWP U10022 ( .A1(n6552), .A2(n6553), .A3(n6554), .A4(n6555), .ZN(
        vectorData2[117]) );
  AOI22D1BWP U10023 ( .A1(n3569), .A2(\vrf/regTable[5][117] ), .B1(n3592), 
        .B2(\vrf/regTable[7][117] ), .ZN(n6555) );
  AOI22D1BWP U10024 ( .A1(n3577), .A2(\vrf/regTable[4][117] ), .B1(n3591), 
        .B2(\vrf/regTable[6][117] ), .ZN(n6554) );
  AOI22D1BWP U10025 ( .A1(n3571), .A2(\vrf/regTable[1][117] ), .B1(n3568), 
        .B2(\vrf/regTable[3][117] ), .ZN(n6553) );
  AOI22D1BWP U10026 ( .A1(n3580), .A2(\vrf/regTable[0][117] ), .B1(n3566), 
        .B2(\vrf/regTable[2][117] ), .ZN(n6552) );
  AOI22D1BWP U10027 ( .A1(n5980), .A2(vectorData2[245]), .B1(n5976), .B2(
        vectorData2[101]), .ZN(n5934) );
  ND4D1BWP U10028 ( .A1(n6488), .A2(n6489), .A3(n6490), .A4(n6491), .ZN(
        vectorData2[101]) );
  AOI22D1BWP U10029 ( .A1(n6082), .A2(\vrf/regTable[5][101] ), .B1(n3578), 
        .B2(\vrf/regTable[7][101] ), .ZN(n6491) );
  AOI22D1BWP U10030 ( .A1(n6080), .A2(\vrf/regTable[4][101] ), .B1(n3573), 
        .B2(\vrf/regTable[6][101] ), .ZN(n6490) );
  AOI22D1BWP U10031 ( .A1(n6077), .A2(\vrf/regTable[1][101] ), .B1(n3597), 
        .B2(\vrf/regTable[3][101] ), .ZN(n6489) );
  AOI22D1BWP U10032 ( .A1(n6073), .A2(\vrf/regTable[0][101] ), .B1(n3593), 
        .B2(\vrf/regTable[2][101] ), .ZN(n6488) );
  ND4D1BWP U10033 ( .A1(n7064), .A2(n7065), .A3(n7066), .A4(n7067), .ZN(
        vectorData2[245]) );
  AOI22D1BWP U10034 ( .A1(n3569), .A2(\vrf/regTable[5][245] ), .B1(n3578), 
        .B2(\vrf/regTable[7][245] ), .ZN(n7067) );
  AOI22D1BWP U10035 ( .A1(n8210), .A2(\vrf/regTable[4][245] ), .B1(n3573), 
        .B2(\vrf/regTable[6][245] ), .ZN(n7066) );
  AOI22D1BWP U10036 ( .A1(n3571), .A2(\vrf/regTable[1][245] ), .B1(n3597), 
        .B2(\vrf/regTable[3][245] ), .ZN(n7065) );
  AOI22D1BWP U10037 ( .A1(n8203), .A2(\vrf/regTable[0][245] ), .B1(n3593), 
        .B2(\vrf/regTable[2][245] ), .ZN(n7064) );
  AOI22D1BWP U10038 ( .A1(n5975), .A2(vectorData2[165]), .B1(n5973), .B2(
        vectorData2[69]), .ZN(n5935) );
  ND4D1BWP U10039 ( .A1(n6360), .A2(n6361), .A3(n6362), .A4(n6363), .ZN(
        vectorData2[69]) );
  AOI22D1BWP U10040 ( .A1(n3569), .A2(\vrf/regTable[5][69] ), .B1(n3578), .B2(
        \vrf/regTable[7][69] ), .ZN(n6363) );
  AOI22D1BWP U10041 ( .A1(n6080), .A2(\vrf/regTable[4][69] ), .B1(n3573), .B2(
        \vrf/regTable[6][69] ), .ZN(n6362) );
  AOI22D1BWP U10042 ( .A1(n3571), .A2(\vrf/regTable[1][69] ), .B1(n3597), .B2(
        \vrf/regTable[3][69] ), .ZN(n6361) );
  AOI22D1BWP U10043 ( .A1(n6073), .A2(\vrf/regTable[0][69] ), .B1(n3593), .B2(
        \vrf/regTable[2][69] ), .ZN(n6360) );
  ND4D1BWP U10044 ( .A1(n6744), .A2(n6745), .A3(n6746), .A4(n6747), .ZN(
        vectorData2[165]) );
  AOI22D1BWP U10045 ( .A1(n3569), .A2(\vrf/regTable[5][165] ), .B1(n3592), 
        .B2(\vrf/regTable[7][165] ), .ZN(n6747) );
  AOI22D1BWP U10046 ( .A1(n8210), .A2(\vrf/regTable[4][165] ), .B1(n3591), 
        .B2(\vrf/regTable[6][165] ), .ZN(n6746) );
  AOI22D1BWP U10047 ( .A1(n3571), .A2(\vrf/regTable[1][165] ), .B1(n3568), 
        .B2(\vrf/regTable[3][165] ), .ZN(n6745) );
  AOI22D1BWP U10048 ( .A1(n8203), .A2(\vrf/regTable[0][165] ), .B1(n3566), 
        .B2(\vrf/regTable[2][165] ), .ZN(n6744) );
  AO22D1BWP U10049 ( .A1(n5977), .A2(vectorData2[133]), .B1(n5983), .B2(
        vectorData2[149]), .Z(n5937) );
  ND4D1BWP U10050 ( .A1(n6680), .A2(n6681), .A3(n6682), .A4(n6683), .ZN(
        vectorData2[149]) );
  AOI22D1BWP U10051 ( .A1(n3569), .A2(\vrf/regTable[5][149] ), .B1(n3578), 
        .B2(\vrf/regTable[7][149] ), .ZN(n6683) );
  AOI22D1BWP U10052 ( .A1(n3577), .A2(\vrf/regTable[4][149] ), .B1(n3573), 
        .B2(\vrf/regTable[6][149] ), .ZN(n6682) );
  AOI22D1BWP U10053 ( .A1(n3571), .A2(\vrf/regTable[1][149] ), .B1(n3597), 
        .B2(\vrf/regTable[3][149] ), .ZN(n6681) );
  AOI22D1BWP U10054 ( .A1(n3580), .A2(\vrf/regTable[0][149] ), .B1(n3593), 
        .B2(\vrf/regTable[2][149] ), .ZN(n6680) );
  ND4D1BWP U10055 ( .A1(n6616), .A2(n6617), .A3(n6618), .A4(n6619), .ZN(
        vectorData2[133]) );
  AOI22D1BWP U10056 ( .A1(n3569), .A2(\vrf/regTable[5][133] ), .B1(n3592), 
        .B2(\vrf/regTable[7][133] ), .ZN(n6619) );
  AOI22D1BWP U10057 ( .A1(n6080), .A2(\vrf/regTable[4][133] ), .B1(n3591), 
        .B2(\vrf/regTable[6][133] ), .ZN(n6618) );
  AOI22D1BWP U10058 ( .A1(n3571), .A2(\vrf/regTable[1][133] ), .B1(n3568), 
        .B2(\vrf/regTable[3][133] ), .ZN(n6617) );
  AOI22D1BWP U10059 ( .A1(n6073), .A2(\vrf/regTable[0][133] ), .B1(n3566), 
        .B2(\vrf/regTable[2][133] ), .ZN(n6616) );
  ND4D1BWP U10060 ( .A1(n6424), .A2(n6425), .A3(n6426), .A4(n6427), .ZN(
        vectorData2[85]) );
  AOI22D1BWP U10061 ( .A1(n3569), .A2(\vrf/regTable[5][85] ), .B1(n3592), .B2(
        \vrf/regTable[7][85] ), .ZN(n6427) );
  AOI22D1BWP U10062 ( .A1(n8210), .A2(\vrf/regTable[4][85] ), .B1(n3591), .B2(
        \vrf/regTable[6][85] ), .ZN(n6426) );
  AOI22D1BWP U10063 ( .A1(n3571), .A2(\vrf/regTable[1][85] ), .B1(n3568), .B2(
        \vrf/regTable[3][85] ), .ZN(n6425) );
  AOI22D1BWP U10064 ( .A1(n8203), .A2(\vrf/regTable[0][85] ), .B1(n3566), .B2(
        \vrf/regTable[2][85] ), .ZN(n6424) );
  AOI22D1BWP U10065 ( .A1(n5974), .A2(vectorData2[53]), .B1(n5984), .B2(
        vectorData2[213]), .ZN(n5939) );
  ND4D1BWP U10066 ( .A1(n6936), .A2(n6937), .A3(n6938), .A4(n6939), .ZN(
        vectorData2[213]) );
  AOI22D1BWP U10067 ( .A1(n3569), .A2(\vrf/regTable[5][213] ), .B1(n3578), 
        .B2(\vrf/regTable[7][213] ), .ZN(n6939) );
  AOI22D1BWP U10068 ( .A1(n3577), .A2(\vrf/regTable[4][213] ), .B1(n3573), 
        .B2(\vrf/regTable[6][213] ), .ZN(n6938) );
  AOI22D1BWP U10069 ( .A1(n3571), .A2(\vrf/regTable[1][213] ), .B1(n3597), 
        .B2(\vrf/regTable[3][213] ), .ZN(n6937) );
  AOI22D1BWP U10070 ( .A1(n3580), .A2(\vrf/regTable[0][213] ), .B1(n3593), 
        .B2(\vrf/regTable[2][213] ), .ZN(n6936) );
  ND4D1BWP U10071 ( .A1(n6296), .A2(n6297), .A3(n6298), .A4(n6299), .ZN(
        vectorData2[53]) );
  AOI22D1BWP U10072 ( .A1(n3569), .A2(\vrf/regTable[5][53] ), .B1(n3592), .B2(
        \vrf/regTable[7][53] ), .ZN(n6299) );
  AOI22D1BWP U10073 ( .A1(n3577), .A2(\vrf/regTable[4][53] ), .B1(n3591), .B2(
        \vrf/regTable[6][53] ), .ZN(n6298) );
  AOI22D1BWP U10074 ( .A1(n3571), .A2(\vrf/regTable[1][53] ), .B1(n3568), .B2(
        \vrf/regTable[3][53] ), .ZN(n6297) );
  AOI22D1BWP U10075 ( .A1(n3580), .A2(\vrf/regTable[0][53] ), .B1(n3566), .B2(
        \vrf/regTable[2][53] ), .ZN(n6296) );
  AOI22D1BWP U10076 ( .A1(n5981), .A2(vectorData2[181]), .B1(n5985), .B2(
        vectorData2[37]), .ZN(n5940) );
  ND4D1BWP U10077 ( .A1(n6232), .A2(n6233), .A3(n6234), .A4(n6235), .ZN(
        vectorData2[37]) );
  AOI22D1BWP U10078 ( .A1(n3569), .A2(\vrf/regTable[5][37] ), .B1(n3578), .B2(
        \vrf/regTable[7][37] ), .ZN(n6235) );
  AOI22D1BWP U10079 ( .A1(n6080), .A2(\vrf/regTable[4][37] ), .B1(n3573), .B2(
        \vrf/regTable[6][37] ), .ZN(n6234) );
  AOI22D1BWP U10080 ( .A1(n3571), .A2(\vrf/regTable[1][37] ), .B1(n3597), .B2(
        \vrf/regTable[3][37] ), .ZN(n6233) );
  AOI22D1BWP U10081 ( .A1(n6073), .A2(\vrf/regTable[0][37] ), .B1(n3593), .B2(
        \vrf/regTable[2][37] ), .ZN(n6232) );
  ND4D1BWP U10082 ( .A1(n6808), .A2(n6809), .A3(n6810), .A4(n6811), .ZN(
        vectorData2[181]) );
  AOI22D1BWP U10083 ( .A1(n3569), .A2(\vrf/regTable[5][181] ), .B1(n3578), 
        .B2(\vrf/regTable[7][181] ), .ZN(n6811) );
  AOI22D1BWP U10084 ( .A1(n3577), .A2(\vrf/regTable[4][181] ), .B1(n3573), 
        .B2(\vrf/regTable[6][181] ), .ZN(n6810) );
  AOI22D1BWP U10085 ( .A1(n3571), .A2(\vrf/regTable[1][181] ), .B1(n3597), 
        .B2(\vrf/regTable[3][181] ), .ZN(n6809) );
  AOI22D1BWP U10086 ( .A1(n3580), .A2(\vrf/regTable[0][181] ), .B1(n3593), 
        .B2(\vrf/regTable[2][181] ), .ZN(n6808) );
  ND4D1BWP U10087 ( .A1(n6104), .A2(n6105), .A3(n6106), .A4(n6107), .ZN(
        vectorData2[5]) );
  AOI22D1BWP U10088 ( .A1(n3569), .A2(\vrf/regTable[5][5] ), .B1(n3592), .B2(
        \vrf/regTable[7][5] ), .ZN(n6107) );
  AOI22D1BWP U10089 ( .A1(n3577), .A2(\vrf/regTable[4][5] ), .B1(n3591), .B2(
        \vrf/regTable[6][5] ), .ZN(n6106) );
  AOI22D1BWP U10090 ( .A1(n3571), .A2(\vrf/regTable[1][5] ), .B1(n3568), .B2(
        \vrf/regTable[3][5] ), .ZN(n6105) );
  AOI22D1BWP U10091 ( .A1(n3580), .A2(\vrf/regTable[0][5] ), .B1(n3566), .B2(
        \vrf/regTable[2][5] ), .ZN(n6104) );
  AO222D1BWP U10092 ( .A1(vectorData2[0]), .A2(n4570), .B1(WR), .B2(n5831), 
        .C1(n4569), .C2(scalarData2[0]), .Z(dataOut[0]) );
  ND4D1BWP U10093 ( .A1(n8214), .A2(n8215), .A3(n8216), .A4(n8217), .ZN(
        scalarData2[0]) );
  AOI22D1BWP U10094 ( .A1(n8212), .A2(\srf/regTable[5][0] ), .B1(n8213), .B2(
        \srf/regTable[7][0] ), .ZN(n8217) );
  AOI22D1BWP U10095 ( .A1(n8210), .A2(\srf/regTable[4][0] ), .B1(n8211), .B2(
        \srf/regTable[6][0] ), .ZN(n8216) );
  AOI22D1BWP U10096 ( .A1(n8207), .A2(\srf/regTable[1][0] ), .B1(n8209), .B2(
        \srf/regTable[3][0] ), .ZN(n8215) );
  AOI22D1BWP U10097 ( .A1(n8203), .A2(\srf/regTable[0][0] ), .B1(n8205), .B2(
        \srf/regTable[2][0] ), .ZN(n8214) );
  ND3D1BWP U10098 ( .A1(n5827), .A2(n5826), .A3(n5825), .ZN(n5831) );
  AOI211XD0BWP U10099 ( .A1(n5981), .A2(vectorData2[176]), .B(n5824), .C(n5823), .ZN(n5825) );
  ND4D1BWP U10100 ( .A1(n5822), .A2(n5821), .A3(n5820), .A4(n5819), .ZN(n5823)
         );
  AOI22D1BWP U10101 ( .A1(n5983), .A2(vectorData2[144]), .B1(n5982), .B2(
        vectorData2[16]), .ZN(n5819) );
  ND4D1BWP U10102 ( .A1(n6148), .A2(n6149), .A3(n6150), .A4(n6151), .ZN(
        vectorData2[16]) );
  AOI22D1BWP U10103 ( .A1(n3569), .A2(\vrf/regTable[5][16] ), .B1(n3592), .B2(
        \vrf/regTable[7][16] ), .ZN(n6151) );
  AOI22D1BWP U10104 ( .A1(n3577), .A2(\vrf/regTable[4][16] ), .B1(n3591), .B2(
        \vrf/regTable[6][16] ), .ZN(n6150) );
  AOI22D1BWP U10105 ( .A1(n3571), .A2(\vrf/regTable[1][16] ), .B1(n3568), .B2(
        \vrf/regTable[3][16] ), .ZN(n6149) );
  AOI22D1BWP U10106 ( .A1(n3580), .A2(\vrf/regTable[0][16] ), .B1(n3566), .B2(
        \vrf/regTable[2][16] ), .ZN(n6148) );
  ND4D1BWP U10107 ( .A1(n6660), .A2(n6661), .A3(n6662), .A4(n6663), .ZN(
        vectorData2[144]) );
  AOI22D1BWP U10108 ( .A1(n3569), .A2(\vrf/regTable[5][144] ), .B1(n3578), 
        .B2(\vrf/regTable[7][144] ), .ZN(n6663) );
  AOI22D1BWP U10109 ( .A1(n3577), .A2(\vrf/regTable[4][144] ), .B1(n3573), 
        .B2(\vrf/regTable[6][144] ), .ZN(n6662) );
  AOI22D1BWP U10110 ( .A1(n3571), .A2(\vrf/regTable[1][144] ), .B1(n3597), 
        .B2(\vrf/regTable[3][144] ), .ZN(n6661) );
  AOI22D1BWP U10111 ( .A1(n3580), .A2(\vrf/regTable[0][144] ), .B1(n3593), 
        .B2(\vrf/regTable[2][144] ), .ZN(n6660) );
  AOI22D1BWP U10112 ( .A1(n5980), .A2(vectorData2[240]), .B1(n5976), .B2(
        vectorData2[96]), .ZN(n5820) );
  ND4D1BWP U10113 ( .A1(n6468), .A2(n6469), .A3(n6470), .A4(n6471), .ZN(
        vectorData2[96]) );
  AOI22D1BWP U10114 ( .A1(n3569), .A2(\vrf/regTable[5][96] ), .B1(n3592), .B2(
        \vrf/regTable[7][96] ), .ZN(n6471) );
  AOI22D1BWP U10115 ( .A1(n6080), .A2(\vrf/regTable[4][96] ), .B1(n3591), .B2(
        \vrf/regTable[6][96] ), .ZN(n6470) );
  AOI22D1BWP U10116 ( .A1(n3571), .A2(\vrf/regTable[1][96] ), .B1(n3568), .B2(
        \vrf/regTable[3][96] ), .ZN(n6469) );
  AOI22D1BWP U10117 ( .A1(n6073), .A2(\vrf/regTable[0][96] ), .B1(n3566), .B2(
        \vrf/regTable[2][96] ), .ZN(n6468) );
  ND4D1BWP U10118 ( .A1(n7044), .A2(n7045), .A3(n7046), .A4(n7047), .ZN(
        vectorData2[240]) );
  AOI22D1BWP U10119 ( .A1(n3569), .A2(\vrf/regTable[5][240] ), .B1(n3592), 
        .B2(\vrf/regTable[7][240] ), .ZN(n7047) );
  AOI22D1BWP U10120 ( .A1(n8210), .A2(\vrf/regTable[4][240] ), .B1(n3591), 
        .B2(\vrf/regTable[6][240] ), .ZN(n7046) );
  AOI22D1BWP U10121 ( .A1(n3571), .A2(\vrf/regTable[1][240] ), .B1(n3568), 
        .B2(\vrf/regTable[3][240] ), .ZN(n7045) );
  AOI22D1BWP U10122 ( .A1(n8203), .A2(\vrf/regTable[0][240] ), .B1(n3566), 
        .B2(\vrf/regTable[2][240] ), .ZN(n7044) );
  AOI22D1BWP U10123 ( .A1(n5978), .A2(vectorData2[192]), .B1(n5973), .B2(
        vectorData2[64]), .ZN(n5821) );
  ND4D1BWP U10124 ( .A1(n6340), .A2(n6341), .A3(n6342), .A4(n6343), .ZN(
        vectorData2[64]) );
  AOI22D1BWP U10125 ( .A1(n3569), .A2(\vrf/regTable[5][64] ), .B1(n3578), .B2(
        \vrf/regTable[7][64] ), .ZN(n6343) );
  AOI22D1BWP U10126 ( .A1(n3577), .A2(\vrf/regTable[4][64] ), .B1(n3573), .B2(
        \vrf/regTable[6][64] ), .ZN(n6342) );
  AOI22D1BWP U10127 ( .A1(n3571), .A2(\vrf/regTable[1][64] ), .B1(n3597), .B2(
        \vrf/regTable[3][64] ), .ZN(n6341) );
  AOI22D1BWP U10128 ( .A1(n3580), .A2(\vrf/regTable[0][64] ), .B1(n3593), .B2(
        \vrf/regTable[2][64] ), .ZN(n6340) );
  ND4D1BWP U10129 ( .A1(n6852), .A2(n6853), .A3(n6854), .A4(n6855), .ZN(
        vectorData2[192]) );
  AOI22D1BWP U10130 ( .A1(n3569), .A2(\vrf/regTable[5][192] ), .B1(n3578), 
        .B2(\vrf/regTable[7][192] ), .ZN(n6855) );
  AOI22D1BWP U10131 ( .A1(n3577), .A2(\vrf/regTable[4][192] ), .B1(n3573), 
        .B2(\vrf/regTable[6][192] ), .ZN(n6854) );
  AOI22D1BWP U10132 ( .A1(n3571), .A2(\vrf/regTable[1][192] ), .B1(n3597), 
        .B2(\vrf/regTable[3][192] ), .ZN(n6853) );
  AOI22D1BWP U10133 ( .A1(n3580), .A2(\vrf/regTable[0][192] ), .B1(n3593), 
        .B2(\vrf/regTable[2][192] ), .ZN(n6852) );
  AOI22D1BWP U10134 ( .A1(n5984), .A2(vectorData2[208]), .B1(n5972), .B2(
        vectorData2[112]), .ZN(n5822) );
  ND4D1BWP U10135 ( .A1(n6532), .A2(n6533), .A3(n6534), .A4(n6535), .ZN(
        vectorData2[112]) );
  AOI22D1BWP U10136 ( .A1(n3569), .A2(\vrf/regTable[5][112] ), .B1(n3578), 
        .B2(\vrf/regTable[7][112] ), .ZN(n6535) );
  AOI22D1BWP U10137 ( .A1(n3577), .A2(\vrf/regTable[4][112] ), .B1(n3573), 
        .B2(\vrf/regTable[6][112] ), .ZN(n6534) );
  AOI22D1BWP U10138 ( .A1(n3571), .A2(\vrf/regTable[1][112] ), .B1(n3597), 
        .B2(\vrf/regTable[3][112] ), .ZN(n6533) );
  AOI22D1BWP U10139 ( .A1(n3580), .A2(\vrf/regTable[0][112] ), .B1(n3593), 
        .B2(\vrf/regTable[2][112] ), .ZN(n6532) );
  ND4D1BWP U10140 ( .A1(n6916), .A2(n6917), .A3(n6918), .A4(n6919), .ZN(
        vectorData2[208]) );
  AOI22D1BWP U10141 ( .A1(n3569), .A2(\vrf/regTable[5][208] ), .B1(n3592), 
        .B2(\vrf/regTable[7][208] ), .ZN(n6919) );
  AOI22D1BWP U10142 ( .A1(n3577), .A2(\vrf/regTable[4][208] ), .B1(n3591), 
        .B2(\vrf/regTable[6][208] ), .ZN(n6918) );
  AOI22D1BWP U10143 ( .A1(n3571), .A2(\vrf/regTable[1][208] ), .B1(n3568), 
        .B2(\vrf/regTable[3][208] ), .ZN(n6917) );
  AOI22D1BWP U10144 ( .A1(n3580), .A2(\vrf/regTable[0][208] ), .B1(n3566), 
        .B2(\vrf/regTable[2][208] ), .ZN(n6916) );
  AO22D1BWP U10145 ( .A1(n5985), .A2(vectorData2[32]), .B1(n5979), .B2(
        vectorData2[80]), .Z(n5824) );
  ND4D1BWP U10146 ( .A1(n6404), .A2(n6405), .A3(n6406), .A4(n6407), .ZN(
        vectorData2[80]) );
  AOI22D1BWP U10147 ( .A1(n3569), .A2(\vrf/regTable[5][80] ), .B1(n3592), .B2(
        \vrf/regTable[7][80] ), .ZN(n6407) );
  AOI22D1BWP U10148 ( .A1(n6080), .A2(\vrf/regTable[4][80] ), .B1(n3591), .B2(
        \vrf/regTable[6][80] ), .ZN(n6406) );
  AOI22D1BWP U10149 ( .A1(n3571), .A2(\vrf/regTable[1][80] ), .B1(n3568), .B2(
        \vrf/regTable[3][80] ), .ZN(n6405) );
  AOI22D1BWP U10150 ( .A1(n6073), .A2(\vrf/regTable[0][80] ), .B1(n3566), .B2(
        \vrf/regTable[2][80] ), .ZN(n6404) );
  ND4D1BWP U10151 ( .A1(n6212), .A2(n6213), .A3(n6214), .A4(n6215), .ZN(
        vectorData2[32]) );
  AOI22D1BWP U10152 ( .A1(n3569), .A2(\vrf/regTable[5][32] ), .B1(n3578), .B2(
        \vrf/regTable[7][32] ), .ZN(n6215) );
  AOI22D1BWP U10153 ( .A1(n3577), .A2(\vrf/regTable[4][32] ), .B1(n3573), .B2(
        \vrf/regTable[6][32] ), .ZN(n6214) );
  AOI22D1BWP U10154 ( .A1(n3571), .A2(\vrf/regTable[1][32] ), .B1(n3597), .B2(
        \vrf/regTable[3][32] ), .ZN(n6213) );
  AOI22D1BWP U10155 ( .A1(n3580), .A2(\vrf/regTable[0][32] ), .B1(n3593), .B2(
        \vrf/regTable[2][32] ), .ZN(n6212) );
  ND4D1BWP U10156 ( .A1(n6788), .A2(n6789), .A3(n6790), .A4(n6791), .ZN(
        vectorData2[176]) );
  AOI22D1BWP U10157 ( .A1(n3569), .A2(\vrf/regTable[5][176] ), .B1(n3578), 
        .B2(\vrf/regTable[7][176] ), .ZN(n6791) );
  AOI22D1BWP U10158 ( .A1(n3577), .A2(\vrf/regTable[4][176] ), .B1(n3573), 
        .B2(\vrf/regTable[6][176] ), .ZN(n6790) );
  AOI22D1BWP U10159 ( .A1(n3571), .A2(\vrf/regTable[1][176] ), .B1(n3597), 
        .B2(\vrf/regTable[3][176] ), .ZN(n6789) );
  AOI22D1BWP U10160 ( .A1(n3580), .A2(\vrf/regTable[0][176] ), .B1(n3593), 
        .B2(\vrf/regTable[2][176] ), .ZN(n6788) );
  AOI22D1BWP U10161 ( .A1(n5992), .A2(vectorData2[224]), .B1(n5975), .B2(
        vectorData2[160]), .ZN(n5826) );
  ND4D1BWP U10162 ( .A1(n6724), .A2(n6725), .A3(n6726), .A4(n6727), .ZN(
        vectorData2[160]) );
  AOI22D1BWP U10163 ( .A1(n3569), .A2(\vrf/regTable[5][160] ), .B1(n3578), 
        .B2(\vrf/regTable[7][160] ), .ZN(n6727) );
  AOI22D1BWP U10164 ( .A1(n3577), .A2(\vrf/regTable[4][160] ), .B1(n3573), 
        .B2(\vrf/regTable[6][160] ), .ZN(n6726) );
  AOI22D1BWP U10165 ( .A1(n3571), .A2(\vrf/regTable[1][160] ), .B1(n3597), 
        .B2(\vrf/regTable[3][160] ), .ZN(n6725) );
  AOI22D1BWP U10166 ( .A1(n3580), .A2(\vrf/regTable[0][160] ), .B1(n3593), 
        .B2(\vrf/regTable[2][160] ), .ZN(n6724) );
  ND4D1BWP U10167 ( .A1(n6980), .A2(n6981), .A3(n6982), .A4(n6983), .ZN(
        vectorData2[224]) );
  AOI22D1BWP U10168 ( .A1(n3569), .A2(\vrf/regTable[5][224] ), .B1(n3592), 
        .B2(\vrf/regTable[7][224] ), .ZN(n6983) );
  AOI22D1BWP U10169 ( .A1(n3577), .A2(\vrf/regTable[4][224] ), .B1(n3591), 
        .B2(\vrf/regTable[6][224] ), .ZN(n6982) );
  AOI22D1BWP U10170 ( .A1(n3571), .A2(\vrf/regTable[1][224] ), .B1(n3568), 
        .B2(\vrf/regTable[3][224] ), .ZN(n6981) );
  AOI22D1BWP U10171 ( .A1(n3580), .A2(\vrf/regTable[0][224] ), .B1(n3566), 
        .B2(\vrf/regTable[2][224] ), .ZN(n6980) );
  AOI22D1BWP U10172 ( .A1(n5974), .A2(vectorData2[48]), .B1(n5977), .B2(
        vectorData2[128]), .ZN(n5827) );
  ND4D1BWP U10173 ( .A1(n6596), .A2(n6597), .A3(n6598), .A4(n6599), .ZN(
        vectorData2[128]) );
  AOI22D1BWP U10174 ( .A1(n3569), .A2(\vrf/regTable[5][128] ), .B1(n3592), 
        .B2(\vrf/regTable[7][128] ), .ZN(n6599) );
  AOI22D1BWP U10175 ( .A1(n8210), .A2(\vrf/regTable[4][128] ), .B1(n3591), 
        .B2(\vrf/regTable[6][128] ), .ZN(n6598) );
  AOI22D1BWP U10176 ( .A1(n3571), .A2(\vrf/regTable[1][128] ), .B1(n3568), 
        .B2(\vrf/regTable[3][128] ), .ZN(n6597) );
  AOI22D1BWP U10177 ( .A1(n8203), .A2(\vrf/regTable[0][128] ), .B1(n3566), 
        .B2(\vrf/regTable[2][128] ), .ZN(n6596) );
  ND4D1BWP U10178 ( .A1(n6276), .A2(n6277), .A3(n6278), .A4(n6279), .ZN(
        vectorData2[48]) );
  AOI22D1BWP U10179 ( .A1(n3569), .A2(\vrf/regTable[5][48] ), .B1(n3578), .B2(
        \vrf/regTable[7][48] ), .ZN(n6279) );
  AOI22D1BWP U10180 ( .A1(n3577), .A2(\vrf/regTable[4][48] ), .B1(n3573), .B2(
        \vrf/regTable[6][48] ), .ZN(n6278) );
  AOI22D1BWP U10181 ( .A1(n3571), .A2(\vrf/regTable[1][48] ), .B1(n3597), .B2(
        \vrf/regTable[3][48] ), .ZN(n6277) );
  AOI22D1BWP U10182 ( .A1(n3580), .A2(\vrf/regTable[0][48] ), .B1(n3593), .B2(
        \vrf/regTable[2][48] ), .ZN(n6276) );
  ND4D1BWP U10183 ( .A1(n6084), .A2(n6085), .A3(n6086), .A4(n6087), .ZN(
        vectorData2[0]) );
  AOI22D1BWP U10184 ( .A1(n3569), .A2(\vrf/regTable[5][0] ), .B1(n3578), .B2(
        \vrf/regTable[7][0] ), .ZN(n6087) );
  AOI22D1BWP U10185 ( .A1(n3577), .A2(\vrf/regTable[4][0] ), .B1(n3573), .B2(
        \vrf/regTable[6][0] ), .ZN(n6086) );
  AOI22D1BWP U10186 ( .A1(n3571), .A2(\vrf/regTable[1][0] ), .B1(n3597), .B2(
        \vrf/regTable[3][0] ), .ZN(n6085) );
  AOI22D1BWP U10187 ( .A1(n3580), .A2(\vrf/regTable[0][0] ), .B1(n3593), .B2(
        \vrf/regTable[2][0] ), .ZN(n6084) );
  AO222D1BWP U10188 ( .A1(vectorData2[7]), .A2(n4570), .B1(WR), .B2(n5961), 
        .C1(scalarData2[7]), .C2(n4569), .Z(dataOut[7]) );
  ND4D1BWP U10189 ( .A1(n8242), .A2(n8243), .A3(n8244), .A4(n8245), .ZN(
        scalarData2[7]) );
  AOI22D1BWP U10190 ( .A1(n8212), .A2(\srf/regTable[5][7] ), .B1(n8213), .B2(
        \srf/regTable[7][7] ), .ZN(n8245) );
  AOI22D1BWP U10191 ( .A1(n8210), .A2(\srf/regTable[4][7] ), .B1(n8211), .B2(
        \srf/regTable[6][7] ), .ZN(n8244) );
  AOI22D1BWP U10192 ( .A1(n8207), .A2(\srf/regTable[1][7] ), .B1(n8209), .B2(
        \srf/regTable[3][7] ), .ZN(n8243) );
  AOI22D1BWP U10193 ( .A1(n8203), .A2(\srf/regTable[0][7] ), .B1(n8205), .B2(
        \srf/regTable[2][7] ), .ZN(n8242) );
  ND3D1BWP U10194 ( .A1(n5960), .A2(n5959), .A3(n5958), .ZN(n5961) );
  AOI211XD0BWP U10195 ( .A1(n5981), .A2(vectorData2[183]), .B(n5957), .C(n5956), .ZN(n5958) );
  ND4D1BWP U10196 ( .A1(n5955), .A2(n5954), .A3(n5953), .A4(n5952), .ZN(n5956)
         );
  AOI22D1BWP U10197 ( .A1(n5975), .A2(vectorData2[167]), .B1(n5976), .B2(
        vectorData2[103]), .ZN(n5952) );
  ND4D1BWP U10198 ( .A1(n6496), .A2(n6497), .A3(n6498), .A4(n6499), .ZN(
        vectorData2[103]) );
  AOI22D1BWP U10199 ( .A1(n3569), .A2(\vrf/regTable[5][103] ), .B1(n3578), 
        .B2(\vrf/regTable[7][103] ), .ZN(n6499) );
  AOI22D1BWP U10200 ( .A1(n3577), .A2(\vrf/regTable[4][103] ), .B1(n3573), 
        .B2(\vrf/regTable[6][103] ), .ZN(n6498) );
  AOI22D1BWP U10201 ( .A1(n3571), .A2(\vrf/regTable[1][103] ), .B1(n3597), 
        .B2(\vrf/regTable[3][103] ), .ZN(n6497) );
  AOI22D1BWP U10202 ( .A1(n3580), .A2(\vrf/regTable[0][103] ), .B1(n3593), 
        .B2(\vrf/regTable[2][103] ), .ZN(n6496) );
  ND4D1BWP U10203 ( .A1(n6752), .A2(n6753), .A3(n6754), .A4(n6755), .ZN(
        vectorData2[167]) );
  AOI22D1BWP U10204 ( .A1(n3569), .A2(\vrf/regTable[5][167] ), .B1(n3592), 
        .B2(\vrf/regTable[7][167] ), .ZN(n6755) );
  AOI22D1BWP U10205 ( .A1(n3577), .A2(\vrf/regTable[4][167] ), .B1(n3591), 
        .B2(\vrf/regTable[6][167] ), .ZN(n6754) );
  AOI22D1BWP U10206 ( .A1(n3571), .A2(\vrf/regTable[1][167] ), .B1(n3568), 
        .B2(\vrf/regTable[3][167] ), .ZN(n6753) );
  AOI22D1BWP U10207 ( .A1(n3580), .A2(\vrf/regTable[0][167] ), .B1(n3566), 
        .B2(\vrf/regTable[2][167] ), .ZN(n6752) );
  AOI22D1BWP U10208 ( .A1(n5974), .A2(vectorData2[55]), .B1(n5972), .B2(
        vectorData2[119]), .ZN(n5953) );
  ND4D1BWP U10209 ( .A1(n6560), .A2(n6561), .A3(n6562), .A4(n6563), .ZN(
        vectorData2[119]) );
  AOI22D1BWP U10210 ( .A1(n3569), .A2(\vrf/regTable[5][119] ), .B1(n3592), 
        .B2(\vrf/regTable[7][119] ), .ZN(n6563) );
  AOI22D1BWP U10211 ( .A1(n3577), .A2(\vrf/regTable[4][119] ), .B1(n3591), 
        .B2(\vrf/regTable[6][119] ), .ZN(n6562) );
  AOI22D1BWP U10212 ( .A1(n3571), .A2(\vrf/regTable[1][119] ), .B1(n3568), 
        .B2(\vrf/regTable[3][119] ), .ZN(n6561) );
  AOI22D1BWP U10213 ( .A1(n3580), .A2(\vrf/regTable[0][119] ), .B1(n3566), 
        .B2(\vrf/regTable[2][119] ), .ZN(n6560) );
  ND4D1BWP U10214 ( .A1(n6304), .A2(n6305), .A3(n6306), .A4(n6307), .ZN(
        vectorData2[55]) );
  AOI22D1BWP U10215 ( .A1(n3569), .A2(\vrf/regTable[5][55] ), .B1(n3592), .B2(
        \vrf/regTable[7][55] ), .ZN(n6307) );
  AOI22D1BWP U10216 ( .A1(n6080), .A2(\vrf/regTable[4][55] ), .B1(n3591), .B2(
        \vrf/regTable[6][55] ), .ZN(n6306) );
  AOI22D1BWP U10217 ( .A1(n3571), .A2(\vrf/regTable[1][55] ), .B1(n3568), .B2(
        \vrf/regTable[3][55] ), .ZN(n6305) );
  AOI22D1BWP U10218 ( .A1(n6073), .A2(\vrf/regTable[0][55] ), .B1(n3566), .B2(
        \vrf/regTable[2][55] ), .ZN(n6304) );
  AOI22D1BWP U10219 ( .A1(n5979), .A2(vectorData2[87]), .B1(n5982), .B2(
        vectorData2[23]), .ZN(n5954) );
  ND4D1BWP U10220 ( .A1(n6176), .A2(n6177), .A3(n6178), .A4(n6179), .ZN(
        vectorData2[23]) );
  AOI22D1BWP U10221 ( .A1(n3569), .A2(\vrf/regTable[5][23] ), .B1(n3578), .B2(
        \vrf/regTable[7][23] ), .ZN(n6179) );
  AOI22D1BWP U10222 ( .A1(n3577), .A2(\vrf/regTable[4][23] ), .B1(n3573), .B2(
        \vrf/regTable[6][23] ), .ZN(n6178) );
  AOI22D1BWP U10223 ( .A1(n3571), .A2(\vrf/regTable[1][23] ), .B1(n3597), .B2(
        \vrf/regTable[3][23] ), .ZN(n6177) );
  AOI22D1BWP U10224 ( .A1(n3580), .A2(\vrf/regTable[0][23] ), .B1(n3593), .B2(
        \vrf/regTable[2][23] ), .ZN(n6176) );
  ND4D1BWP U10225 ( .A1(n6432), .A2(n6433), .A3(n6434), .A4(n6435), .ZN(
        vectorData2[87]) );
  AOI22D1BWP U10226 ( .A1(n6082), .A2(\vrf/regTable[5][87] ), .B1(n3592), .B2(
        \vrf/regTable[7][87] ), .ZN(n6435) );
  AOI22D1BWP U10227 ( .A1(n6080), .A2(\vrf/regTable[4][87] ), .B1(n3591), .B2(
        \vrf/regTable[6][87] ), .ZN(n6434) );
  AOI22D1BWP U10228 ( .A1(n6077), .A2(\vrf/regTable[1][87] ), .B1(n3568), .B2(
        \vrf/regTable[3][87] ), .ZN(n6433) );
  AOI22D1BWP U10229 ( .A1(n6073), .A2(\vrf/regTable[0][87] ), .B1(n3566), .B2(
        \vrf/regTable[2][87] ), .ZN(n6432) );
  AOI22D1BWP U10230 ( .A1(n5977), .A2(vectorData2[135]), .B1(n5983), .B2(
        vectorData2[151]), .ZN(n5955) );
  ND4D1BWP U10231 ( .A1(n6688), .A2(n6689), .A3(n6690), .A4(n6691), .ZN(
        vectorData2[151]) );
  AOI22D1BWP U10232 ( .A1(n3569), .A2(\vrf/regTable[5][151] ), .B1(n3578), 
        .B2(\vrf/regTable[7][151] ), .ZN(n6691) );
  AOI22D1BWP U10233 ( .A1(n3577), .A2(\vrf/regTable[4][151] ), .B1(n3573), 
        .B2(\vrf/regTable[6][151] ), .ZN(n6690) );
  AOI22D1BWP U10234 ( .A1(n3571), .A2(\vrf/regTable[1][151] ), .B1(n3597), 
        .B2(\vrf/regTable[3][151] ), .ZN(n6689) );
  AOI22D1BWP U10235 ( .A1(n3580), .A2(\vrf/regTable[0][151] ), .B1(n3593), 
        .B2(\vrf/regTable[2][151] ), .ZN(n6688) );
  ND4D1BWP U10236 ( .A1(n6624), .A2(n6625), .A3(n6626), .A4(n6627), .ZN(
        vectorData2[135]) );
  AOI22D1BWP U10237 ( .A1(n3569), .A2(\vrf/regTable[5][135] ), .B1(n3592), 
        .B2(\vrf/regTable[7][135] ), .ZN(n6627) );
  AOI22D1BWP U10238 ( .A1(n8210), .A2(\vrf/regTable[4][135] ), .B1(n3591), 
        .B2(\vrf/regTable[6][135] ), .ZN(n6626) );
  AOI22D1BWP U10239 ( .A1(n3571), .A2(\vrf/regTable[1][135] ), .B1(n3568), 
        .B2(\vrf/regTable[3][135] ), .ZN(n6625) );
  AOI22D1BWP U10240 ( .A1(n8203), .A2(\vrf/regTable[0][135] ), .B1(n3566), 
        .B2(\vrf/regTable[2][135] ), .ZN(n6624) );
  AO22D1BWP U10241 ( .A1(n5985), .A2(vectorData2[39]), .B1(n5992), .B2(
        vectorData2[231]), .Z(n5957) );
  ND4D1BWP U10242 ( .A1(n7008), .A2(n7009), .A3(n7010), .A4(n7011), .ZN(
        vectorData2[231]) );
  AOI22D1BWP U10243 ( .A1(n3569), .A2(\vrf/regTable[5][231] ), .B1(n3578), 
        .B2(\vrf/regTable[7][231] ), .ZN(n7011) );
  AOI22D1BWP U10244 ( .A1(n3577), .A2(\vrf/regTable[4][231] ), .B1(n3573), 
        .B2(\vrf/regTable[6][231] ), .ZN(n7010) );
  AOI22D1BWP U10245 ( .A1(n3571), .A2(\vrf/regTable[1][231] ), .B1(n3597), 
        .B2(\vrf/regTable[3][231] ), .ZN(n7009) );
  AOI22D1BWP U10246 ( .A1(n3580), .A2(\vrf/regTable[0][231] ), .B1(n3593), 
        .B2(\vrf/regTable[2][231] ), .ZN(n7008) );
  ND4D1BWP U10247 ( .A1(n6240), .A2(n6241), .A3(n6242), .A4(n6243), .ZN(
        vectorData2[39]) );
  AOI22D1BWP U10248 ( .A1(n3569), .A2(\vrf/regTable[5][39] ), .B1(n3592), .B2(
        \vrf/regTable[7][39] ), .ZN(n6243) );
  AOI22D1BWP U10249 ( .A1(n3577), .A2(\vrf/regTable[4][39] ), .B1(n3591), .B2(
        \vrf/regTable[6][39] ), .ZN(n6242) );
  AOI22D1BWP U10250 ( .A1(n3571), .A2(\vrf/regTable[1][39] ), .B1(n3568), .B2(
        \vrf/regTable[3][39] ), .ZN(n6241) );
  AOI22D1BWP U10251 ( .A1(n3580), .A2(\vrf/regTable[0][39] ), .B1(n3566), .B2(
        \vrf/regTable[2][39] ), .ZN(n6240) );
  ND4D1BWP U10252 ( .A1(n6816), .A2(n6817), .A3(n6818), .A4(n6819), .ZN(
        vectorData2[183]) );
  AOI22D1BWP U10253 ( .A1(n3569), .A2(\vrf/regTable[5][183] ), .B1(n3592), 
        .B2(\vrf/regTable[7][183] ), .ZN(n6819) );
  AOI22D1BWP U10254 ( .A1(n3577), .A2(\vrf/regTable[4][183] ), .B1(n3591), 
        .B2(\vrf/regTable[6][183] ), .ZN(n6818) );
  AOI22D1BWP U10255 ( .A1(n3571), .A2(\vrf/regTable[1][183] ), .B1(n3568), 
        .B2(\vrf/regTable[3][183] ), .ZN(n6817) );
  AOI22D1BWP U10256 ( .A1(n3580), .A2(\vrf/regTable[0][183] ), .B1(n3566), 
        .B2(\vrf/regTable[2][183] ), .ZN(n6816) );
  AOI22D1BWP U10257 ( .A1(n5978), .A2(vectorData2[199]), .B1(n5973), .B2(
        vectorData2[71]), .ZN(n5959) );
  ND4D1BWP U10258 ( .A1(n6368), .A2(n6369), .A3(n6370), .A4(n6371), .ZN(
        vectorData2[71]) );
  AOI22D1BWP U10259 ( .A1(n3569), .A2(\vrf/regTable[5][71] ), .B1(n3592), .B2(
        \vrf/regTable[7][71] ), .ZN(n6371) );
  AOI22D1BWP U10260 ( .A1(n3577), .A2(\vrf/regTable[4][71] ), .B1(n3591), .B2(
        \vrf/regTable[6][71] ), .ZN(n6370) );
  AOI22D1BWP U10261 ( .A1(n3571), .A2(\vrf/regTable[1][71] ), .B1(n3568), .B2(
        \vrf/regTable[3][71] ), .ZN(n6369) );
  AOI22D1BWP U10262 ( .A1(n3580), .A2(\vrf/regTable[0][71] ), .B1(n3566), .B2(
        \vrf/regTable[2][71] ), .ZN(n6368) );
  ND4D1BWP U10263 ( .A1(n6880), .A2(n6881), .A3(n6882), .A4(n6883), .ZN(
        vectorData2[199]) );
  AOI22D1BWP U10264 ( .A1(n3569), .A2(\vrf/regTable[5][199] ), .B1(n3592), 
        .B2(\vrf/regTable[7][199] ), .ZN(n6883) );
  AOI22D1BWP U10265 ( .A1(n3577), .A2(\vrf/regTable[4][199] ), .B1(n3591), 
        .B2(\vrf/regTable[6][199] ), .ZN(n6882) );
  AOI22D1BWP U10266 ( .A1(n3571), .A2(\vrf/regTable[1][199] ), .B1(n3568), 
        .B2(\vrf/regTable[3][199] ), .ZN(n6881) );
  AOI22D1BWP U10267 ( .A1(n3580), .A2(\vrf/regTable[0][199] ), .B1(n3566), 
        .B2(\vrf/regTable[2][199] ), .ZN(n6880) );
  AOI22D1BWP U10268 ( .A1(n5984), .A2(vectorData2[215]), .B1(n5980), .B2(
        vectorData2[247]), .ZN(n5960) );
  ND4D1BWP U10269 ( .A1(n7072), .A2(n7073), .A3(n7074), .A4(n7075), .ZN(
        vectorData2[247]) );
  AOI22D1BWP U10270 ( .A1(n3569), .A2(\vrf/regTable[5][247] ), .B1(n6083), 
        .B2(\vrf/regTable[7][247] ), .ZN(n7075) );
  AOI22D1BWP U10271 ( .A1(n3577), .A2(\vrf/regTable[4][247] ), .B1(n6081), 
        .B2(\vrf/regTable[6][247] ), .ZN(n7074) );
  AOI22D1BWP U10272 ( .A1(n3571), .A2(\vrf/regTable[1][247] ), .B1(n6079), 
        .B2(\vrf/regTable[3][247] ), .ZN(n7073) );
  AOI22D1BWP U10273 ( .A1(n3580), .A2(\vrf/regTable[0][247] ), .B1(n6075), 
        .B2(\vrf/regTable[2][247] ), .ZN(n7072) );
  ND4D1BWP U10274 ( .A1(n6944), .A2(n6945), .A3(n6946), .A4(n6947), .ZN(
        vectorData2[215]) );
  AOI22D1BWP U10275 ( .A1(n3569), .A2(\vrf/regTable[5][215] ), .B1(n3578), 
        .B2(\vrf/regTable[7][215] ), .ZN(n6947) );
  AOI22D1BWP U10276 ( .A1(n3577), .A2(\vrf/regTable[4][215] ), .B1(n3573), 
        .B2(\vrf/regTable[6][215] ), .ZN(n6946) );
  AOI22D1BWP U10277 ( .A1(n3571), .A2(\vrf/regTable[1][215] ), .B1(n3597), 
        .B2(\vrf/regTable[3][215] ), .ZN(n6945) );
  AOI22D1BWP U10278 ( .A1(n3580), .A2(\vrf/regTable[0][215] ), .B1(n3593), 
        .B2(\vrf/regTable[2][215] ), .ZN(n6944) );
  ND4D1BWP U10279 ( .A1(n6112), .A2(n6113), .A3(n6114), .A4(n6115), .ZN(
        vectorData2[7]) );
  AOI22D1BWP U10280 ( .A1(n3569), .A2(\vrf/regTable[5][7] ), .B1(n3592), .B2(
        \vrf/regTable[7][7] ), .ZN(n6115) );
  AOI22D1BWP U10281 ( .A1(n3577), .A2(\vrf/regTable[4][7] ), .B1(n3591), .B2(
        \vrf/regTable[6][7] ), .ZN(n6114) );
  AOI22D1BWP U10282 ( .A1(n3571), .A2(\vrf/regTable[1][7] ), .B1(n3568), .B2(
        \vrf/regTable[3][7] ), .ZN(n6113) );
  AOI22D1BWP U10283 ( .A1(n3580), .A2(\vrf/regTable[0][7] ), .B1(n3566), .B2(
        \vrf/regTable[2][7] ), .ZN(n6112) );
  AO222D1BWP U10284 ( .A1(WR), .A2(n5911), .B1(n4570), .B2(vectorData2[2]), 
        .C1(n4569), .C2(scalarData2[2]), .Z(dataOut[2]) );
  ND4D1BWP U10285 ( .A1(n8222), .A2(n8223), .A3(n8224), .A4(n8225), .ZN(
        scalarData2[2]) );
  AOI22D1BWP U10286 ( .A1(n8212), .A2(\srf/regTable[5][2] ), .B1(n8213), .B2(
        \srf/regTable[7][2] ), .ZN(n8225) );
  AOI22D1BWP U10287 ( .A1(n8210), .A2(\srf/regTable[4][2] ), .B1(n8211), .B2(
        \srf/regTable[6][2] ), .ZN(n8224) );
  AOI22D1BWP U10288 ( .A1(n8207), .A2(\srf/regTable[1][2] ), .B1(n8209), .B2(
        \srf/regTable[3][2] ), .ZN(n8223) );
  AOI22D1BWP U10289 ( .A1(n8203), .A2(\srf/regTable[0][2] ), .B1(n8205), .B2(
        \srf/regTable[2][2] ), .ZN(n8222) );
  ND4D1BWP U10290 ( .A1(n6092), .A2(n6093), .A3(n6094), .A4(n6095), .ZN(
        vectorData2[2]) );
  AOI22D1BWP U10291 ( .A1(n3569), .A2(\vrf/regTable[5][2] ), .B1(n3578), .B2(
        \vrf/regTable[7][2] ), .ZN(n6095) );
  AOI22D1BWP U10292 ( .A1(n3577), .A2(\vrf/regTable[4][2] ), .B1(n3573), .B2(
        \vrf/regTable[6][2] ), .ZN(n6094) );
  AOI22D1BWP U10293 ( .A1(n3571), .A2(\vrf/regTable[1][2] ), .B1(n3597), .B2(
        \vrf/regTable[3][2] ), .ZN(n6093) );
  AOI22D1BWP U10294 ( .A1(n3580), .A2(\vrf/regTable[0][2] ), .B1(n3593), .B2(
        \vrf/regTable[2][2] ), .ZN(n6092) );
  ND3D1BWP U10295 ( .A1(n5910), .A2(n5909), .A3(n5908), .ZN(n5911) );
  AOI211XD0BWP U10296 ( .A1(n5974), .A2(vectorData2[50]), .B(n5907), .C(n5906), 
        .ZN(n5908) );
  ND4D1BWP U10297 ( .A1(n5905), .A2(n5904), .A3(n5903), .A4(n5902), .ZN(n5906)
         );
  AOI22D1BWP U10298 ( .A1(n5984), .A2(vectorData2[210]), .B1(n5982), .B2(
        vectorData2[18]), .ZN(n5902) );
  ND4D1BWP U10299 ( .A1(n6156), .A2(n6157), .A3(n6158), .A4(n6159), .ZN(
        vectorData2[18]) );
  AOI22D1BWP U10300 ( .A1(n3569), .A2(\vrf/regTable[5][18] ), .B1(n3592), .B2(
        \vrf/regTable[7][18] ), .ZN(n6159) );
  AOI22D1BWP U10301 ( .A1(n3577), .A2(\vrf/regTable[4][18] ), .B1(n3591), .B2(
        \vrf/regTable[6][18] ), .ZN(n6158) );
  AOI22D1BWP U10302 ( .A1(n3571), .A2(\vrf/regTable[1][18] ), .B1(n3568), .B2(
        \vrf/regTable[3][18] ), .ZN(n6157) );
  AOI22D1BWP U10303 ( .A1(n3580), .A2(\vrf/regTable[0][18] ), .B1(n3566), .B2(
        \vrf/regTable[2][18] ), .ZN(n6156) );
  ND4D1BWP U10304 ( .A1(n6924), .A2(n6925), .A3(n6926), .A4(n6927), .ZN(
        vectorData2[210]) );
  AOI22D1BWP U10305 ( .A1(n3569), .A2(\vrf/regTable[5][210] ), .B1(n6083), 
        .B2(\vrf/regTable[7][210] ), .ZN(n6927) );
  AOI22D1BWP U10306 ( .A1(n3577), .A2(\vrf/regTable[4][210] ), .B1(n6081), 
        .B2(\vrf/regTable[6][210] ), .ZN(n6926) );
  AOI22D1BWP U10307 ( .A1(n3571), .A2(\vrf/regTable[1][210] ), .B1(n6079), 
        .B2(\vrf/regTable[3][210] ), .ZN(n6925) );
  AOI22D1BWP U10308 ( .A1(n3580), .A2(\vrf/regTable[0][210] ), .B1(n6075), 
        .B2(\vrf/regTable[2][210] ), .ZN(n6924) );
  AOI22D1BWP U10309 ( .A1(n5981), .A2(vectorData2[178]), .B1(n5980), .B2(
        vectorData2[242]), .ZN(n5903) );
  ND4D1BWP U10310 ( .A1(n7052), .A2(n7053), .A3(n7054), .A4(n7055), .ZN(
        vectorData2[242]) );
  AOI22D1BWP U10311 ( .A1(n3569), .A2(\vrf/regTable[5][242] ), .B1(n3592), 
        .B2(\vrf/regTable[7][242] ), .ZN(n7055) );
  AOI22D1BWP U10312 ( .A1(n6080), .A2(\vrf/regTable[4][242] ), .B1(n3591), 
        .B2(\vrf/regTable[6][242] ), .ZN(n7054) );
  AOI22D1BWP U10313 ( .A1(n3571), .A2(\vrf/regTable[1][242] ), .B1(n3568), 
        .B2(\vrf/regTable[3][242] ), .ZN(n7053) );
  AOI22D1BWP U10314 ( .A1(n6073), .A2(\vrf/regTable[0][242] ), .B1(n3566), 
        .B2(\vrf/regTable[2][242] ), .ZN(n7052) );
  ND4D1BWP U10315 ( .A1(n6796), .A2(n6797), .A3(n6798), .A4(n6799), .ZN(
        vectorData2[178]) );
  AOI22D1BWP U10316 ( .A1(n3569), .A2(\vrf/regTable[5][178] ), .B1(n3578), 
        .B2(\vrf/regTable[7][178] ), .ZN(n6799) );
  AOI22D1BWP U10317 ( .A1(n3577), .A2(\vrf/regTable[4][178] ), .B1(n3573), 
        .B2(\vrf/regTable[6][178] ), .ZN(n6798) );
  AOI22D1BWP U10318 ( .A1(n3571), .A2(\vrf/regTable[1][178] ), .B1(n3597), 
        .B2(\vrf/regTable[3][178] ), .ZN(n6797) );
  AOI22D1BWP U10319 ( .A1(n3580), .A2(\vrf/regTable[0][178] ), .B1(n3593), 
        .B2(\vrf/regTable[2][178] ), .ZN(n6796) );
  AOI22D1BWP U10320 ( .A1(n5978), .A2(vectorData2[194]), .B1(n5972), .B2(
        vectorData2[114]), .ZN(n5904) );
  ND4D1BWP U10321 ( .A1(n6540), .A2(n6541), .A3(n6542), .A4(n6543), .ZN(
        vectorData2[114]) );
  AOI22D1BWP U10322 ( .A1(n3569), .A2(\vrf/regTable[5][114] ), .B1(n3578), 
        .B2(\vrf/regTable[7][114] ), .ZN(n6543) );
  AOI22D1BWP U10323 ( .A1(n3577), .A2(\vrf/regTable[4][114] ), .B1(n3573), 
        .B2(\vrf/regTable[6][114] ), .ZN(n6542) );
  AOI22D1BWP U10324 ( .A1(n3571), .A2(\vrf/regTable[1][114] ), .B1(n3597), 
        .B2(\vrf/regTable[3][114] ), .ZN(n6541) );
  AOI22D1BWP U10325 ( .A1(n3580), .A2(\vrf/regTable[0][114] ), .B1(n3593), 
        .B2(\vrf/regTable[2][114] ), .ZN(n6540) );
  ND4D1BWP U10326 ( .A1(n6860), .A2(n6861), .A3(n6862), .A4(n6863), .ZN(
        vectorData2[194]) );
  AOI22D1BWP U10327 ( .A1(n3569), .A2(\vrf/regTable[5][194] ), .B1(n3592), 
        .B2(\vrf/regTable[7][194] ), .ZN(n6863) );
  AOI22D1BWP U10328 ( .A1(n3577), .A2(\vrf/regTable[4][194] ), .B1(n3591), 
        .B2(\vrf/regTable[6][194] ), .ZN(n6862) );
  AOI22D1BWP U10329 ( .A1(n3571), .A2(\vrf/regTable[1][194] ), .B1(n3568), 
        .B2(\vrf/regTable[3][194] ), .ZN(n6861) );
  AOI22D1BWP U10330 ( .A1(n3580), .A2(\vrf/regTable[0][194] ), .B1(n3566), 
        .B2(\vrf/regTable[2][194] ), .ZN(n6860) );
  AOI22D1BWP U10331 ( .A1(n5975), .A2(vectorData2[162]), .B1(n5976), .B2(
        vectorData2[98]), .ZN(n5905) );
  ND4D1BWP U10332 ( .A1(n6476), .A2(n6477), .A3(n6478), .A4(n6479), .ZN(
        vectorData2[98]) );
  AOI22D1BWP U10333 ( .A1(n3569), .A2(\vrf/regTable[5][98] ), .B1(n3592), .B2(
        \vrf/regTable[7][98] ), .ZN(n6479) );
  AOI22D1BWP U10334 ( .A1(n3577), .A2(\vrf/regTable[4][98] ), .B1(n3591), .B2(
        \vrf/regTable[6][98] ), .ZN(n6478) );
  AOI22D1BWP U10335 ( .A1(n3571), .A2(\vrf/regTable[1][98] ), .B1(n3568), .B2(
        \vrf/regTable[3][98] ), .ZN(n6477) );
  AOI22D1BWP U10336 ( .A1(n3580), .A2(\vrf/regTable[0][98] ), .B1(n3566), .B2(
        \vrf/regTable[2][98] ), .ZN(n6476) );
  ND4D1BWP U10337 ( .A1(n6732), .A2(n6733), .A3(n6734), .A4(n6735), .ZN(
        vectorData2[162]) );
  AOI22D1BWP U10338 ( .A1(n3569), .A2(\vrf/regTable[5][162] ), .B1(n3592), 
        .B2(\vrf/regTable[7][162] ), .ZN(n6735) );
  AOI22D1BWP U10339 ( .A1(n8210), .A2(\vrf/regTable[4][162] ), .B1(n3591), 
        .B2(\vrf/regTable[6][162] ), .ZN(n6734) );
  AOI22D1BWP U10340 ( .A1(n3571), .A2(\vrf/regTable[1][162] ), .B1(n3568), 
        .B2(\vrf/regTable[3][162] ), .ZN(n6733) );
  AOI22D1BWP U10341 ( .A1(n8203), .A2(\vrf/regTable[0][162] ), .B1(n3566), 
        .B2(\vrf/regTable[2][162] ), .ZN(n6732) );
  AO22D1BWP U10342 ( .A1(n5973), .A2(vectorData2[66]), .B1(n5983), .B2(
        vectorData2[146]), .Z(n5907) );
  ND4D1BWP U10343 ( .A1(n6668), .A2(n6669), .A3(n6670), .A4(n6671), .ZN(
        vectorData2[146]) );
  AOI22D1BWP U10344 ( .A1(n3569), .A2(\vrf/regTable[5][146] ), .B1(n3578), 
        .B2(\vrf/regTable[7][146] ), .ZN(n6671) );
  AOI22D1BWP U10345 ( .A1(n6080), .A2(\vrf/regTable[4][146] ), .B1(n3573), 
        .B2(\vrf/regTable[6][146] ), .ZN(n6670) );
  AOI22D1BWP U10346 ( .A1(n3571), .A2(\vrf/regTable[1][146] ), .B1(n3597), 
        .B2(\vrf/regTable[3][146] ), .ZN(n6669) );
  AOI22D1BWP U10347 ( .A1(n6073), .A2(\vrf/regTable[0][146] ), .B1(n3593), 
        .B2(\vrf/regTable[2][146] ), .ZN(n6668) );
  ND4D1BWP U10348 ( .A1(n6348), .A2(n6349), .A3(n6350), .A4(n6351), .ZN(
        vectorData2[66]) );
  AOI22D1BWP U10349 ( .A1(n6082), .A2(\vrf/regTable[5][66] ), .B1(n3592), .B2(
        \vrf/regTable[7][66] ), .ZN(n6351) );
  AOI22D1BWP U10350 ( .A1(n6080), .A2(\vrf/regTable[4][66] ), .B1(n3591), .B2(
        \vrf/regTable[6][66] ), .ZN(n6350) );
  AOI22D1BWP U10351 ( .A1(n6077), .A2(\vrf/regTable[1][66] ), .B1(n3568), .B2(
        \vrf/regTable[3][66] ), .ZN(n6349) );
  AOI22D1BWP U10352 ( .A1(n6073), .A2(\vrf/regTable[0][66] ), .B1(n3566), .B2(
        \vrf/regTable[2][66] ), .ZN(n6348) );
  ND4D1BWP U10353 ( .A1(n6284), .A2(n6285), .A3(n6286), .A4(n6287), .ZN(
        vectorData2[50]) );
  AOI22D1BWP U10354 ( .A1(n3569), .A2(\vrf/regTable[5][50] ), .B1(n3578), .B2(
        \vrf/regTable[7][50] ), .ZN(n6287) );
  AOI22D1BWP U10355 ( .A1(n3577), .A2(\vrf/regTable[4][50] ), .B1(n3573), .B2(
        \vrf/regTable[6][50] ), .ZN(n6286) );
  AOI22D1BWP U10356 ( .A1(n3571), .A2(\vrf/regTable[1][50] ), .B1(n3597), .B2(
        \vrf/regTable[3][50] ), .ZN(n6285) );
  AOI22D1BWP U10357 ( .A1(n3580), .A2(\vrf/regTable[0][50] ), .B1(n3593), .B2(
        \vrf/regTable[2][50] ), .ZN(n6284) );
  AOI22D1BWP U10358 ( .A1(n5985), .A2(vectorData2[34]), .B1(n5992), .B2(
        vectorData2[226]), .ZN(n5909) );
  ND4D1BWP U10359 ( .A1(n6988), .A2(n6989), .A3(n6990), .A4(n6991), .ZN(
        vectorData2[226]) );
  AOI22D1BWP U10360 ( .A1(n3569), .A2(\vrf/regTable[5][226] ), .B1(n3592), 
        .B2(\vrf/regTable[7][226] ), .ZN(n6991) );
  AOI22D1BWP U10361 ( .A1(n8210), .A2(\vrf/regTable[4][226] ), .B1(n3591), 
        .B2(\vrf/regTable[6][226] ), .ZN(n6990) );
  AOI22D1BWP U10362 ( .A1(n3571), .A2(\vrf/regTable[1][226] ), .B1(n3568), 
        .B2(\vrf/regTable[3][226] ), .ZN(n6989) );
  AOI22D1BWP U10363 ( .A1(n8203), .A2(\vrf/regTable[0][226] ), .B1(n3566), 
        .B2(\vrf/regTable[2][226] ), .ZN(n6988) );
  ND4D1BWP U10364 ( .A1(n6220), .A2(n6221), .A3(n6222), .A4(n6223), .ZN(
        vectorData2[34]) );
  AOI22D1BWP U10365 ( .A1(n3569), .A2(\vrf/regTable[5][34] ), .B1(n3578), .B2(
        \vrf/regTable[7][34] ), .ZN(n6223) );
  AOI22D1BWP U10366 ( .A1(n3577), .A2(\vrf/regTable[4][34] ), .B1(n3573), .B2(
        \vrf/regTable[6][34] ), .ZN(n6222) );
  AOI22D1BWP U10367 ( .A1(n3571), .A2(\vrf/regTable[1][34] ), .B1(n3597), .B2(
        \vrf/regTable[3][34] ), .ZN(n6221) );
  AOI22D1BWP U10368 ( .A1(n3580), .A2(\vrf/regTable[0][34] ), .B1(n3593), .B2(
        \vrf/regTable[2][34] ), .ZN(n6220) );
  AOI22D1BWP U10369 ( .A1(n5979), .A2(vectorData2[82]), .B1(n5977), .B2(
        vectorData2[130]), .ZN(n5910) );
  ND4D1BWP U10370 ( .A1(n6604), .A2(n6605), .A3(n6606), .A4(n6607), .ZN(
        vectorData2[130]) );
  AOI22D1BWP U10371 ( .A1(n3569), .A2(\vrf/regTable[5][130] ), .B1(n3592), 
        .B2(\vrf/regTable[7][130] ), .ZN(n6607) );
  AOI22D1BWP U10372 ( .A1(n3577), .A2(\vrf/regTable[4][130] ), .B1(n3591), 
        .B2(\vrf/regTable[6][130] ), .ZN(n6606) );
  AOI22D1BWP U10373 ( .A1(n3571), .A2(\vrf/regTable[1][130] ), .B1(n3568), 
        .B2(\vrf/regTable[3][130] ), .ZN(n6605) );
  AOI22D1BWP U10374 ( .A1(n3580), .A2(\vrf/regTable[0][130] ), .B1(n3566), 
        .B2(\vrf/regTable[2][130] ), .ZN(n6604) );
  ND4D1BWP U10375 ( .A1(n6412), .A2(n6413), .A3(n6414), .A4(n6415), .ZN(
        vectorData2[82]) );
  AOI22D1BWP U10376 ( .A1(n6082), .A2(\vrf/regTable[5][82] ), .B1(n3592), .B2(
        \vrf/regTable[7][82] ), .ZN(n6415) );
  AOI22D1BWP U10377 ( .A1(n6080), .A2(\vrf/regTable[4][82] ), .B1(n3591), .B2(
        \vrf/regTable[6][82] ), .ZN(n6414) );
  AOI22D1BWP U10378 ( .A1(n6077), .A2(\vrf/regTable[1][82] ), .B1(n3568), .B2(
        \vrf/regTable[3][82] ), .ZN(n6413) );
  AOI22D1BWP U10379 ( .A1(n6073), .A2(\vrf/regTable[0][82] ), .B1(n3566), .B2(
        \vrf/regTable[2][82] ), .ZN(n6412) );
  AO222D1BWP U10380 ( .A1(vectorData2[3]), .A2(n4570), .B1(WR), .B2(n5921), 
        .C1(scalarData2[3]), .C2(n4569), .Z(dataOut[3]) );
  ND4D1BWP U10381 ( .A1(n8226), .A2(n8227), .A3(n8228), .A4(n8229), .ZN(
        scalarData2[3]) );
  AOI22D1BWP U10382 ( .A1(n8212), .A2(\srf/regTable[5][3] ), .B1(n8213), .B2(
        \srf/regTable[7][3] ), .ZN(n8229) );
  AOI22D1BWP U10383 ( .A1(n8210), .A2(\srf/regTable[4][3] ), .B1(n8211), .B2(
        \srf/regTable[6][3] ), .ZN(n8228) );
  AOI22D1BWP U10384 ( .A1(n8207), .A2(\srf/regTable[1][3] ), .B1(n8209), .B2(
        \srf/regTable[3][3] ), .ZN(n8227) );
  AOI22D1BWP U10385 ( .A1(n8203), .A2(\srf/regTable[0][3] ), .B1(n8205), .B2(
        \srf/regTable[2][3] ), .ZN(n8226) );
  ND3D1BWP U10386 ( .A1(n5920), .A2(n5919), .A3(n5918), .ZN(n5921) );
  AOI211XD0BWP U10387 ( .A1(n5979), .A2(vectorData2[83]), .B(n5917), .C(n5916), 
        .ZN(n5918) );
  ND4D1BWP U10388 ( .A1(n5915), .A2(n5914), .A3(n5913), .A4(n5912), .ZN(n5916)
         );
  AOI22D1BWP U10389 ( .A1(n5973), .A2(vectorData2[67]), .B1(n5984), .B2(
        vectorData2[211]), .ZN(n5912) );
  ND4D1BWP U10390 ( .A1(n6928), .A2(n6929), .A3(n6930), .A4(n6931), .ZN(
        vectorData2[211]) );
  AOI22D1BWP U10391 ( .A1(n3569), .A2(\vrf/regTable[5][211] ), .B1(n6083), 
        .B2(\vrf/regTable[7][211] ), .ZN(n6931) );
  AOI22D1BWP U10392 ( .A1(n3577), .A2(\vrf/regTable[4][211] ), .B1(n6081), 
        .B2(\vrf/regTable[6][211] ), .ZN(n6930) );
  AOI22D1BWP U10393 ( .A1(n3571), .A2(\vrf/regTable[1][211] ), .B1(n6079), 
        .B2(\vrf/regTable[3][211] ), .ZN(n6929) );
  AOI22D1BWP U10394 ( .A1(n3580), .A2(\vrf/regTable[0][211] ), .B1(n6075), 
        .B2(\vrf/regTable[2][211] ), .ZN(n6928) );
  ND4D1BWP U10395 ( .A1(n6352), .A2(n6353), .A3(n6354), .A4(n6355), .ZN(
        vectorData2[67]) );
  AOI22D1BWP U10396 ( .A1(n3569), .A2(\vrf/regTable[5][67] ), .B1(n3578), .B2(
        \vrf/regTable[7][67] ), .ZN(n6355) );
  AOI22D1BWP U10397 ( .A1(n3577), .A2(\vrf/regTable[4][67] ), .B1(n3573), .B2(
        \vrf/regTable[6][67] ), .ZN(n6354) );
  AOI22D1BWP U10398 ( .A1(n3571), .A2(\vrf/regTable[1][67] ), .B1(n3597), .B2(
        \vrf/regTable[3][67] ), .ZN(n6353) );
  AOI22D1BWP U10399 ( .A1(n3580), .A2(\vrf/regTable[0][67] ), .B1(n3593), .B2(
        \vrf/regTable[2][67] ), .ZN(n6352) );
  AOI22D1BWP U10400 ( .A1(n5985), .A2(vectorData2[35]), .B1(n5992), .B2(
        vectorData2[227]), .ZN(n5913) );
  ND4D1BWP U10401 ( .A1(n6992), .A2(n6993), .A3(n6994), .A4(n6995), .ZN(
        vectorData2[227]) );
  AOI22D1BWP U10402 ( .A1(n3569), .A2(\vrf/regTable[5][227] ), .B1(n3592), 
        .B2(\vrf/regTable[7][227] ), .ZN(n6995) );
  AOI22D1BWP U10403 ( .A1(n3577), .A2(\vrf/regTable[4][227] ), .B1(n3591), 
        .B2(\vrf/regTable[6][227] ), .ZN(n6994) );
  AOI22D1BWP U10404 ( .A1(n3571), .A2(\vrf/regTable[1][227] ), .B1(n3568), 
        .B2(\vrf/regTable[3][227] ), .ZN(n6993) );
  AOI22D1BWP U10405 ( .A1(n3580), .A2(\vrf/regTable[0][227] ), .B1(n3566), 
        .B2(\vrf/regTable[2][227] ), .ZN(n6992) );
  ND4D1BWP U10406 ( .A1(n6224), .A2(n6225), .A3(n6226), .A4(n6227), .ZN(
        vectorData2[35]) );
  AOI22D1BWP U10407 ( .A1(n3569), .A2(\vrf/regTable[5][35] ), .B1(n3592), .B2(
        \vrf/regTable[7][35] ), .ZN(n6227) );
  AOI22D1BWP U10408 ( .A1(n3577), .A2(\vrf/regTable[4][35] ), .B1(n3591), .B2(
        \vrf/regTable[6][35] ), .ZN(n6226) );
  AOI22D1BWP U10409 ( .A1(n3571), .A2(\vrf/regTable[1][35] ), .B1(n3568), .B2(
        \vrf/regTable[3][35] ), .ZN(n6225) );
  AOI22D1BWP U10410 ( .A1(n3580), .A2(\vrf/regTable[0][35] ), .B1(n3566), .B2(
        \vrf/regTable[2][35] ), .ZN(n6224) );
  AOI22D1BWP U10411 ( .A1(n5981), .A2(vectorData2[179]), .B1(n5977), .B2(
        vectorData2[131]), .ZN(n5914) );
  ND4D1BWP U10412 ( .A1(n6608), .A2(n6609), .A3(n6610), .A4(n6611), .ZN(
        vectorData2[131]) );
  AOI22D1BWP U10413 ( .A1(n3569), .A2(\vrf/regTable[5][131] ), .B1(n3592), 
        .B2(\vrf/regTable[7][131] ), .ZN(n6611) );
  AOI22D1BWP U10414 ( .A1(n3577), .A2(\vrf/regTable[4][131] ), .B1(n3591), 
        .B2(\vrf/regTable[6][131] ), .ZN(n6610) );
  AOI22D1BWP U10415 ( .A1(n3571), .A2(\vrf/regTable[1][131] ), .B1(n3568), 
        .B2(\vrf/regTable[3][131] ), .ZN(n6609) );
  AOI22D1BWP U10416 ( .A1(n3580), .A2(\vrf/regTable[0][131] ), .B1(n3566), 
        .B2(\vrf/regTable[2][131] ), .ZN(n6608) );
  ND4D1BWP U10417 ( .A1(n6800), .A2(n6801), .A3(n6802), .A4(n6803), .ZN(
        vectorData2[179]) );
  AOI22D1BWP U10418 ( .A1(n3569), .A2(\vrf/regTable[5][179] ), .B1(n3578), 
        .B2(\vrf/regTable[7][179] ), .ZN(n6803) );
  AOI22D1BWP U10419 ( .A1(n3577), .A2(\vrf/regTable[4][179] ), .B1(n3573), 
        .B2(\vrf/regTable[6][179] ), .ZN(n6802) );
  AOI22D1BWP U10420 ( .A1(n3571), .A2(\vrf/regTable[1][179] ), .B1(n3597), 
        .B2(\vrf/regTable[3][179] ), .ZN(n6801) );
  AOI22D1BWP U10421 ( .A1(n3580), .A2(\vrf/regTable[0][179] ), .B1(n3593), 
        .B2(\vrf/regTable[2][179] ), .ZN(n6800) );
  AOI22D1BWP U10422 ( .A1(n5972), .A2(vectorData2[115]), .B1(n5980), .B2(
        vectorData2[243]), .ZN(n5915) );
  ND4D1BWP U10423 ( .A1(n7056), .A2(n7057), .A3(n7058), .A4(n7059), .ZN(
        vectorData2[243]) );
  AOI22D1BWP U10424 ( .A1(n3569), .A2(\vrf/regTable[5][243] ), .B1(n3592), 
        .B2(\vrf/regTable[7][243] ), .ZN(n7059) );
  AOI22D1BWP U10425 ( .A1(n6080), .A2(\vrf/regTable[4][243] ), .B1(n3591), 
        .B2(\vrf/regTable[6][243] ), .ZN(n7058) );
  AOI22D1BWP U10426 ( .A1(n3571), .A2(\vrf/regTable[1][243] ), .B1(n3568), 
        .B2(\vrf/regTable[3][243] ), .ZN(n7057) );
  AOI22D1BWP U10427 ( .A1(n6073), .A2(\vrf/regTable[0][243] ), .B1(n3566), 
        .B2(\vrf/regTable[2][243] ), .ZN(n7056) );
  ND4D1BWP U10428 ( .A1(n6544), .A2(n6545), .A3(n6546), .A4(n6547), .ZN(
        vectorData2[115]) );
  AOI22D1BWP U10429 ( .A1(n3569), .A2(\vrf/regTable[5][115] ), .B1(n3592), 
        .B2(\vrf/regTable[7][115] ), .ZN(n6547) );
  AOI22D1BWP U10430 ( .A1(n3577), .A2(\vrf/regTable[4][115] ), .B1(n3591), 
        .B2(\vrf/regTable[6][115] ), .ZN(n6546) );
  AOI22D1BWP U10431 ( .A1(n3571), .A2(\vrf/regTable[1][115] ), .B1(n3568), 
        .B2(\vrf/regTable[3][115] ), .ZN(n6545) );
  AOI22D1BWP U10432 ( .A1(n3580), .A2(\vrf/regTable[0][115] ), .B1(n3566), 
        .B2(\vrf/regTable[2][115] ), .ZN(n6544) );
  AO22D1BWP U10433 ( .A1(n5975), .A2(vectorData2[163]), .B1(n5982), .B2(
        vectorData2[19]), .Z(n5917) );
  ND4D1BWP U10434 ( .A1(n6160), .A2(n6161), .A3(n6162), .A4(n6163), .ZN(
        vectorData2[19]) );
  AOI22D1BWP U10435 ( .A1(n6082), .A2(\vrf/regTable[5][19] ), .B1(n3578), .B2(
        \vrf/regTable[7][19] ), .ZN(n6163) );
  AOI22D1BWP U10436 ( .A1(n3577), .A2(\vrf/regTable[4][19] ), .B1(n3573), .B2(
        \vrf/regTable[6][19] ), .ZN(n6162) );
  AOI22D1BWP U10437 ( .A1(n6077), .A2(\vrf/regTable[1][19] ), .B1(n3597), .B2(
        \vrf/regTable[3][19] ), .ZN(n6161) );
  AOI22D1BWP U10438 ( .A1(n3580), .A2(\vrf/regTable[0][19] ), .B1(n3593), .B2(
        \vrf/regTable[2][19] ), .ZN(n6160) );
  ND4D1BWP U10439 ( .A1(n6736), .A2(n6737), .A3(n6738), .A4(n6739), .ZN(
        vectorData2[163]) );
  AOI22D1BWP U10440 ( .A1(n3569), .A2(\vrf/regTable[5][163] ), .B1(n3578), 
        .B2(\vrf/regTable[7][163] ), .ZN(n6739) );
  AOI22D1BWP U10441 ( .A1(n3577), .A2(\vrf/regTable[4][163] ), .B1(n3573), 
        .B2(\vrf/regTable[6][163] ), .ZN(n6738) );
  AOI22D1BWP U10442 ( .A1(n3571), .A2(\vrf/regTable[1][163] ), .B1(n3597), 
        .B2(\vrf/regTable[3][163] ), .ZN(n6737) );
  AOI22D1BWP U10443 ( .A1(n3580), .A2(\vrf/regTable[0][163] ), .B1(n3593), 
        .B2(\vrf/regTable[2][163] ), .ZN(n6736) );
  ND4D1BWP U10444 ( .A1(n6416), .A2(n6417), .A3(n6418), .A4(n6419), .ZN(
        vectorData2[83]) );
  AOI22D1BWP U10445 ( .A1(n3569), .A2(\vrf/regTable[5][83] ), .B1(n3578), .B2(
        \vrf/regTable[7][83] ), .ZN(n6419) );
  AOI22D1BWP U10446 ( .A1(n3577), .A2(\vrf/regTable[4][83] ), .B1(n3573), .B2(
        \vrf/regTable[6][83] ), .ZN(n6418) );
  AOI22D1BWP U10447 ( .A1(n3571), .A2(\vrf/regTable[1][83] ), .B1(n3597), .B2(
        \vrf/regTable[3][83] ), .ZN(n6417) );
  AOI22D1BWP U10448 ( .A1(n3580), .A2(\vrf/regTable[0][83] ), .B1(n3593), .B2(
        \vrf/regTable[2][83] ), .ZN(n6416) );
  AOI22D1BWP U10449 ( .A1(n5974), .A2(vectorData2[51]), .B1(n5983), .B2(
        vectorData2[147]), .ZN(n5919) );
  ND4D1BWP U10450 ( .A1(n6672), .A2(n6673), .A3(n6674), .A4(n6675), .ZN(
        vectorData2[147]) );
  AOI22D1BWP U10451 ( .A1(n3569), .A2(\vrf/regTable[5][147] ), .B1(n3578), 
        .B2(\vrf/regTable[7][147] ), .ZN(n6675) );
  AOI22D1BWP U10452 ( .A1(n3577), .A2(\vrf/regTable[4][147] ), .B1(n3573), 
        .B2(\vrf/regTable[6][147] ), .ZN(n6674) );
  AOI22D1BWP U10453 ( .A1(n3571), .A2(\vrf/regTable[1][147] ), .B1(n3597), 
        .B2(\vrf/regTable[3][147] ), .ZN(n6673) );
  AOI22D1BWP U10454 ( .A1(n3580), .A2(\vrf/regTable[0][147] ), .B1(n3593), 
        .B2(\vrf/regTable[2][147] ), .ZN(n6672) );
  ND4D1BWP U10455 ( .A1(n6288), .A2(n6289), .A3(n6290), .A4(n6291), .ZN(
        vectorData2[51]) );
  AOI22D1BWP U10456 ( .A1(n3569), .A2(\vrf/regTable[5][51] ), .B1(n3578), .B2(
        \vrf/regTable[7][51] ), .ZN(n6291) );
  AOI22D1BWP U10457 ( .A1(n3577), .A2(\vrf/regTable[4][51] ), .B1(n3573), .B2(
        \vrf/regTable[6][51] ), .ZN(n6290) );
  AOI22D1BWP U10458 ( .A1(n3571), .A2(\vrf/regTable[1][51] ), .B1(n3597), .B2(
        \vrf/regTable[3][51] ), .ZN(n6289) );
  AOI22D1BWP U10459 ( .A1(n3580), .A2(\vrf/regTable[0][51] ), .B1(n3593), .B2(
        \vrf/regTable[2][51] ), .ZN(n6288) );
  AOI22D1BWP U10460 ( .A1(n5978), .A2(vectorData2[195]), .B1(n5976), .B2(
        vectorData2[99]), .ZN(n5920) );
  ND4D1BWP U10461 ( .A1(n6480), .A2(n6481), .A3(n6482), .A4(n6483), .ZN(
        vectorData2[99]) );
  AOI22D1BWP U10462 ( .A1(n3569), .A2(\vrf/regTable[5][99] ), .B1(n3592), .B2(
        \vrf/regTable[7][99] ), .ZN(n6483) );
  AOI22D1BWP U10463 ( .A1(n3577), .A2(\vrf/regTable[4][99] ), .B1(n3591), .B2(
        \vrf/regTable[6][99] ), .ZN(n6482) );
  AOI22D1BWP U10464 ( .A1(n3571), .A2(\vrf/regTable[1][99] ), .B1(n3568), .B2(
        \vrf/regTable[3][99] ), .ZN(n6481) );
  AOI22D1BWP U10465 ( .A1(n3580), .A2(\vrf/regTable[0][99] ), .B1(n3566), .B2(
        \vrf/regTable[2][99] ), .ZN(n6480) );
  ND4D1BWP U10466 ( .A1(n6864), .A2(n6865), .A3(n6866), .A4(n6867), .ZN(
        vectorData2[195]) );
  AOI22D1BWP U10467 ( .A1(n3569), .A2(\vrf/regTable[5][195] ), .B1(n3578), 
        .B2(\vrf/regTable[7][195] ), .ZN(n6867) );
  AOI22D1BWP U10468 ( .A1(n3577), .A2(\vrf/regTable[4][195] ), .B1(n3573), 
        .B2(\vrf/regTable[6][195] ), .ZN(n6866) );
  AOI22D1BWP U10469 ( .A1(n3571), .A2(\vrf/regTable[1][195] ), .B1(n3597), 
        .B2(\vrf/regTable[3][195] ), .ZN(n6865) );
  AOI22D1BWP U10470 ( .A1(n3580), .A2(\vrf/regTable[0][195] ), .B1(n3593), 
        .B2(\vrf/regTable[2][195] ), .ZN(n6864) );
  ND4D1BWP U10471 ( .A1(n6096), .A2(n6097), .A3(n6098), .A4(n6099), .ZN(
        vectorData2[3]) );
  AOI22D1BWP U10472 ( .A1(n3569), .A2(\vrf/regTable[5][3] ), .B1(n3578), .B2(
        \vrf/regTable[7][3] ), .ZN(n6099) );
  AOI22D1BWP U10473 ( .A1(n3577), .A2(\vrf/regTable[4][3] ), .B1(n3573), .B2(
        \vrf/regTable[6][3] ), .ZN(n6098) );
  AOI22D1BWP U10474 ( .A1(n3571), .A2(\vrf/regTable[1][3] ), .B1(n3597), .B2(
        \vrf/regTable[3][3] ), .ZN(n6097) );
  AOI22D1BWP U10475 ( .A1(n3580), .A2(\vrf/regTable[0][3] ), .B1(n3593), .B2(
        \vrf/regTable[2][3] ), .ZN(n6096) );
  AO222D1BWP U10476 ( .A1(WR), .A2(n5861), .B1(n4570), .B2(vectorData2[12]), 
        .C1(n4569), .C2(scalarData2[12]), .Z(dataOut[12]) );
  ND4D1BWP U10477 ( .A1(n8262), .A2(n8263), .A3(n8264), .A4(n8265), .ZN(
        scalarData2[12]) );
  AOI22D1BWP U10478 ( .A1(n8212), .A2(\srf/regTable[5][12] ), .B1(n8213), .B2(
        \srf/regTable[7][12] ), .ZN(n8265) );
  AOI22D1BWP U10479 ( .A1(n8210), .A2(\srf/regTable[4][12] ), .B1(n8211), .B2(
        \srf/regTable[6][12] ), .ZN(n8264) );
  AOI22D1BWP U10480 ( .A1(n8207), .A2(\srf/regTable[1][12] ), .B1(n8209), .B2(
        \srf/regTable[3][12] ), .ZN(n8263) );
  AOI22D1BWP U10481 ( .A1(n8203), .A2(\srf/regTable[0][12] ), .B1(n8205), .B2(
        \srf/regTable[2][12] ), .ZN(n8262) );
  ND4D1BWP U10482 ( .A1(n6132), .A2(n6133), .A3(n6134), .A4(n6135), .ZN(
        vectorData2[12]) );
  AOI22D1BWP U10483 ( .A1(n3569), .A2(\vrf/regTable[5][12] ), .B1(n3578), .B2(
        \vrf/regTable[7][12] ), .ZN(n6135) );
  AOI22D1BWP U10484 ( .A1(n8210), .A2(\vrf/regTable[4][12] ), .B1(n3573), .B2(
        \vrf/regTable[6][12] ), .ZN(n6134) );
  AOI22D1BWP U10485 ( .A1(n3571), .A2(\vrf/regTable[1][12] ), .B1(n3597), .B2(
        \vrf/regTable[3][12] ), .ZN(n6133) );
  AOI22D1BWP U10486 ( .A1(n8203), .A2(\vrf/regTable[0][12] ), .B1(n3593), .B2(
        \vrf/regTable[2][12] ), .ZN(n6132) );
  ND3D1BWP U10487 ( .A1(n5860), .A2(n5859), .A3(n5858), .ZN(n5861) );
  AOI211XD0BWP U10488 ( .A1(n5978), .A2(vectorData2[204]), .B(n5857), .C(n5856), .ZN(n5858) );
  ND4D1BWP U10489 ( .A1(n5855), .A2(n5854), .A3(n5853), .A4(n5852), .ZN(n5856)
         );
  AOI22D1BWP U10490 ( .A1(n5985), .A2(vectorData2[44]), .B1(n5979), .B2(
        vectorData2[92]), .ZN(n5852) );
  ND4D1BWP U10491 ( .A1(n6452), .A2(n6453), .A3(n6454), .A4(n6455), .ZN(
        vectorData2[92]) );
  AOI22D1BWP U10492 ( .A1(n6082), .A2(\vrf/regTable[5][92] ), .B1(n3592), .B2(
        \vrf/regTable[7][92] ), .ZN(n6455) );
  AOI22D1BWP U10493 ( .A1(n6080), .A2(\vrf/regTable[4][92] ), .B1(n3591), .B2(
        \vrf/regTable[6][92] ), .ZN(n6454) );
  AOI22D1BWP U10494 ( .A1(n6077), .A2(\vrf/regTable[1][92] ), .B1(n3568), .B2(
        \vrf/regTable[3][92] ), .ZN(n6453) );
  AOI22D1BWP U10495 ( .A1(n6073), .A2(\vrf/regTable[0][92] ), .B1(n3566), .B2(
        \vrf/regTable[2][92] ), .ZN(n6452) );
  ND4D1BWP U10496 ( .A1(n6260), .A2(n6261), .A3(n6262), .A4(n6263), .ZN(
        vectorData2[44]) );
  AOI22D1BWP U10497 ( .A1(n3569), .A2(\vrf/regTable[5][44] ), .B1(n3578), .B2(
        \vrf/regTable[7][44] ), .ZN(n6263) );
  AOI22D1BWP U10498 ( .A1(n6080), .A2(\vrf/regTable[4][44] ), .B1(n3573), .B2(
        \vrf/regTable[6][44] ), .ZN(n6262) );
  AOI22D1BWP U10499 ( .A1(n3571), .A2(\vrf/regTable[1][44] ), .B1(n3597), .B2(
        \vrf/regTable[3][44] ), .ZN(n6261) );
  AOI22D1BWP U10500 ( .A1(n6073), .A2(\vrf/regTable[0][44] ), .B1(n3593), .B2(
        \vrf/regTable[2][44] ), .ZN(n6260) );
  AOI22D1BWP U10501 ( .A1(n5974), .A2(vectorData2[60]), .B1(n5983), .B2(
        vectorData2[156]), .ZN(n5853) );
  ND4D1BWP U10502 ( .A1(n6708), .A2(n6709), .A3(n6710), .A4(n6711), .ZN(
        vectorData2[156]) );
  AOI22D1BWP U10503 ( .A1(n3569), .A2(\vrf/regTable[5][156] ), .B1(n3592), 
        .B2(\vrf/regTable[7][156] ), .ZN(n6711) );
  AOI22D1BWP U10504 ( .A1(n6080), .A2(\vrf/regTable[4][156] ), .B1(n3591), 
        .B2(\vrf/regTable[6][156] ), .ZN(n6710) );
  AOI22D1BWP U10505 ( .A1(n3571), .A2(\vrf/regTable[1][156] ), .B1(n3568), 
        .B2(\vrf/regTable[3][156] ), .ZN(n6709) );
  AOI22D1BWP U10506 ( .A1(n6073), .A2(\vrf/regTable[0][156] ), .B1(n3566), 
        .B2(\vrf/regTable[2][156] ), .ZN(n6708) );
  ND4D1BWP U10507 ( .A1(n6324), .A2(n6325), .A3(n6326), .A4(n6327), .ZN(
        vectorData2[60]) );
  AOI22D1BWP U10508 ( .A1(n3569), .A2(\vrf/regTable[5][60] ), .B1(n3592), .B2(
        \vrf/regTable[7][60] ), .ZN(n6327) );
  AOI22D1BWP U10509 ( .A1(n8210), .A2(\vrf/regTable[4][60] ), .B1(n3591), .B2(
        \vrf/regTable[6][60] ), .ZN(n6326) );
  AOI22D1BWP U10510 ( .A1(n3571), .A2(\vrf/regTable[1][60] ), .B1(n3568), .B2(
        \vrf/regTable[3][60] ), .ZN(n6325) );
  AOI22D1BWP U10511 ( .A1(n8203), .A2(\vrf/regTable[0][60] ), .B1(n3566), .B2(
        \vrf/regTable[2][60] ), .ZN(n6324) );
  AOI22D1BWP U10512 ( .A1(n5992), .A2(vectorData2[236]), .B1(n5973), .B2(
        vectorData2[76]), .ZN(n5854) );
  ND4D1BWP U10513 ( .A1(n6388), .A2(n6389), .A3(n6390), .A4(n6391), .ZN(
        vectorData2[76]) );
  AOI22D1BWP U10514 ( .A1(n3569), .A2(\vrf/regTable[5][76] ), .B1(n3592), .B2(
        \vrf/regTable[7][76] ), .ZN(n6391) );
  AOI22D1BWP U10515 ( .A1(n3577), .A2(\vrf/regTable[4][76] ), .B1(n3591), .B2(
        \vrf/regTable[6][76] ), .ZN(n6390) );
  AOI22D1BWP U10516 ( .A1(n3571), .A2(\vrf/regTable[1][76] ), .B1(n3568), .B2(
        \vrf/regTable[3][76] ), .ZN(n6389) );
  AOI22D1BWP U10517 ( .A1(n3580), .A2(\vrf/regTable[0][76] ), .B1(n3566), .B2(
        \vrf/regTable[2][76] ), .ZN(n6388) );
  ND4D1BWP U10518 ( .A1(n7028), .A2(n7029), .A3(n7030), .A4(n7031), .ZN(
        vectorData2[236]) );
  AOI22D1BWP U10519 ( .A1(n3569), .A2(\vrf/regTable[5][236] ), .B1(n3578), 
        .B2(\vrf/regTable[7][236] ), .ZN(n7031) );
  AOI22D1BWP U10520 ( .A1(n6080), .A2(\vrf/regTable[4][236] ), .B1(n3573), 
        .B2(\vrf/regTable[6][236] ), .ZN(n7030) );
  AOI22D1BWP U10521 ( .A1(n3571), .A2(\vrf/regTable[1][236] ), .B1(n3597), 
        .B2(\vrf/regTable[3][236] ), .ZN(n7029) );
  AOI22D1BWP U10522 ( .A1(n6073), .A2(\vrf/regTable[0][236] ), .B1(n3593), 
        .B2(\vrf/regTable[2][236] ), .ZN(n7028) );
  AOI22D1BWP U10523 ( .A1(n5977), .A2(vectorData2[140]), .B1(n5972), .B2(
        vectorData2[124]), .ZN(n5855) );
  ND4D1BWP U10524 ( .A1(n6580), .A2(n6581), .A3(n6582), .A4(n6583), .ZN(
        vectorData2[124]) );
  AOI22D1BWP U10525 ( .A1(n6082), .A2(\vrf/regTable[5][124] ), .B1(n3592), 
        .B2(\vrf/regTable[7][124] ), .ZN(n6583) );
  AOI22D1BWP U10526 ( .A1(n6080), .A2(\vrf/regTable[4][124] ), .B1(n3591), 
        .B2(\vrf/regTable[6][124] ), .ZN(n6582) );
  AOI22D1BWP U10527 ( .A1(n6077), .A2(\vrf/regTable[1][124] ), .B1(n3568), 
        .B2(\vrf/regTable[3][124] ), .ZN(n6581) );
  AOI22D1BWP U10528 ( .A1(n6073), .A2(\vrf/regTable[0][124] ), .B1(n3566), 
        .B2(\vrf/regTable[2][124] ), .ZN(n6580) );
  ND4D1BWP U10529 ( .A1(n6644), .A2(n6645), .A3(n6646), .A4(n6647), .ZN(
        vectorData2[140]) );
  AOI22D1BWP U10530 ( .A1(n3569), .A2(\vrf/regTable[5][140] ), .B1(n3592), 
        .B2(\vrf/regTable[7][140] ), .ZN(n6647) );
  AOI22D1BWP U10531 ( .A1(n3577), .A2(\vrf/regTable[4][140] ), .B1(n3591), 
        .B2(\vrf/regTable[6][140] ), .ZN(n6646) );
  AOI22D1BWP U10532 ( .A1(n3571), .A2(\vrf/regTable[1][140] ), .B1(n3568), 
        .B2(\vrf/regTable[3][140] ), .ZN(n6645) );
  AOI22D1BWP U10533 ( .A1(n3580), .A2(\vrf/regTable[0][140] ), .B1(n3566), 
        .B2(\vrf/regTable[2][140] ), .ZN(n6644) );
  AO22D1BWP U10534 ( .A1(n5980), .A2(vectorData2[252]), .B1(n5976), .B2(
        vectorData2[108]), .Z(n5857) );
  ND4D1BWP U10535 ( .A1(n6516), .A2(n6517), .A3(n6518), .A4(n6519), .ZN(
        vectorData2[108]) );
  AOI22D1BWP U10536 ( .A1(n3569), .A2(\vrf/regTable[5][108] ), .B1(n3578), 
        .B2(\vrf/regTable[7][108] ), .ZN(n6519) );
  AOI22D1BWP U10537 ( .A1(n3577), .A2(\vrf/regTable[4][108] ), .B1(n3573), 
        .B2(\vrf/regTable[6][108] ), .ZN(n6518) );
  AOI22D1BWP U10538 ( .A1(n3571), .A2(\vrf/regTable[1][108] ), .B1(n3597), 
        .B2(\vrf/regTable[3][108] ), .ZN(n6517) );
  AOI22D1BWP U10539 ( .A1(n3580), .A2(\vrf/regTable[0][108] ), .B1(n3593), 
        .B2(\vrf/regTable[2][108] ), .ZN(n6516) );
  ND4D1BWP U10540 ( .A1(n7092), .A2(n7093), .A3(n7094), .A4(n7095), .ZN(
        vectorData2[252]) );
  AOI22D1BWP U10541 ( .A1(n3569), .A2(\vrf/regTable[5][252] ), .B1(n6083), 
        .B2(\vrf/regTable[7][252] ), .ZN(n7095) );
  AOI22D1BWP U10542 ( .A1(n8210), .A2(\vrf/regTable[4][252] ), .B1(n6081), 
        .B2(\vrf/regTable[6][252] ), .ZN(n7094) );
  AOI22D1BWP U10543 ( .A1(n3571), .A2(\vrf/regTable[1][252] ), .B1(n6079), 
        .B2(\vrf/regTable[3][252] ), .ZN(n7093) );
  AOI22D1BWP U10544 ( .A1(n8203), .A2(\vrf/regTable[0][252] ), .B1(n6075), 
        .B2(\vrf/regTable[2][252] ), .ZN(n7092) );
  ND4D1BWP U10545 ( .A1(n6900), .A2(n6901), .A3(n6902), .A4(n6903), .ZN(
        vectorData2[204]) );
  AOI22D1BWP U10546 ( .A1(n3569), .A2(\vrf/regTable[5][204] ), .B1(n6083), 
        .B2(\vrf/regTable[7][204] ), .ZN(n6903) );
  AOI22D1BWP U10547 ( .A1(n3577), .A2(\vrf/regTable[4][204] ), .B1(n6081), 
        .B2(\vrf/regTable[6][204] ), .ZN(n6902) );
  AOI22D1BWP U10548 ( .A1(n3571), .A2(\vrf/regTable[1][204] ), .B1(n6079), 
        .B2(\vrf/regTable[3][204] ), .ZN(n6901) );
  AOI22D1BWP U10549 ( .A1(n3580), .A2(\vrf/regTable[0][204] ), .B1(n6075), 
        .B2(\vrf/regTable[2][204] ), .ZN(n6900) );
  AOI22D1BWP U10550 ( .A1(n5981), .A2(vectorData2[188]), .B1(n5984), .B2(
        vectorData2[220]), .ZN(n5859) );
  ND4D1BWP U10551 ( .A1(n6964), .A2(n6965), .A3(n6966), .A4(n6967), .ZN(
        vectorData2[220]) );
  AOI22D1BWP U10552 ( .A1(n3569), .A2(\vrf/regTable[5][220] ), .B1(n6083), 
        .B2(\vrf/regTable[7][220] ), .ZN(n6967) );
  AOI22D1BWP U10553 ( .A1(n6080), .A2(\vrf/regTable[4][220] ), .B1(n6081), 
        .B2(\vrf/regTable[6][220] ), .ZN(n6966) );
  AOI22D1BWP U10554 ( .A1(n3571), .A2(\vrf/regTable[1][220] ), .B1(n6079), 
        .B2(\vrf/regTable[3][220] ), .ZN(n6965) );
  AOI22D1BWP U10555 ( .A1(n6073), .A2(\vrf/regTable[0][220] ), .B1(n6075), 
        .B2(\vrf/regTable[2][220] ), .ZN(n6964) );
  ND4D1BWP U10556 ( .A1(n6836), .A2(n6837), .A3(n6838), .A4(n6839), .ZN(
        vectorData2[188]) );
  AOI22D1BWP U10557 ( .A1(n3569), .A2(\vrf/regTable[5][188] ), .B1(n3592), 
        .B2(\vrf/regTable[7][188] ), .ZN(n6839) );
  AOI22D1BWP U10558 ( .A1(n3577), .A2(\vrf/regTable[4][188] ), .B1(n3591), 
        .B2(\vrf/regTable[6][188] ), .ZN(n6838) );
  AOI22D1BWP U10559 ( .A1(n3571), .A2(\vrf/regTable[1][188] ), .B1(n3568), 
        .B2(\vrf/regTable[3][188] ), .ZN(n6837) );
  AOI22D1BWP U10560 ( .A1(n3580), .A2(\vrf/regTable[0][188] ), .B1(n3566), 
        .B2(\vrf/regTable[2][188] ), .ZN(n6836) );
  AOI22D1BWP U10561 ( .A1(n5975), .A2(vectorData2[172]), .B1(n5982), .B2(
        vectorData2[28]), .ZN(n5860) );
  ND4D1BWP U10562 ( .A1(n6196), .A2(n6197), .A3(n6198), .A4(n6199), .ZN(
        vectorData2[28]) );
  AOI22D1BWP U10563 ( .A1(n3569), .A2(\vrf/regTable[5][28] ), .B1(n3578), .B2(
        \vrf/regTable[7][28] ), .ZN(n6199) );
  AOI22D1BWP U10564 ( .A1(n3577), .A2(\vrf/regTable[4][28] ), .B1(n3573), .B2(
        \vrf/regTable[6][28] ), .ZN(n6198) );
  AOI22D1BWP U10565 ( .A1(n3571), .A2(\vrf/regTable[1][28] ), .B1(n3597), .B2(
        \vrf/regTable[3][28] ), .ZN(n6197) );
  AOI22D1BWP U10566 ( .A1(n3580), .A2(\vrf/regTable[0][28] ), .B1(n3593), .B2(
        \vrf/regTable[2][28] ), .ZN(n6196) );
  ND4D1BWP U10567 ( .A1(n6772), .A2(n6773), .A3(n6774), .A4(n6775), .ZN(
        vectorData2[172]) );
  AOI22D1BWP U10568 ( .A1(n3569), .A2(\vrf/regTable[5][172] ), .B1(n3578), 
        .B2(\vrf/regTable[7][172] ), .ZN(n6775) );
  AOI22D1BWP U10569 ( .A1(n3577), .A2(\vrf/regTable[4][172] ), .B1(n3573), 
        .B2(\vrf/regTable[6][172] ), .ZN(n6774) );
  AOI22D1BWP U10570 ( .A1(n3571), .A2(\vrf/regTable[1][172] ), .B1(n3597), 
        .B2(\vrf/regTable[3][172] ), .ZN(n6773) );
  AOI22D1BWP U10571 ( .A1(n3580), .A2(\vrf/regTable[0][172] ), .B1(n3593), 
        .B2(\vrf/regTable[2][172] ), .ZN(n6772) );
  AO222D1BWP U10572 ( .A1(WR), .A2(n5871), .B1(n4570), .B2(vectorData2[13]), 
        .C1(n4569), .C2(scalarData2[13]), .Z(dataOut[13]) );
  ND4D1BWP U10573 ( .A1(n8266), .A2(n8267), .A3(n8268), .A4(n8269), .ZN(
        scalarData2[13]) );
  AOI22D1BWP U10574 ( .A1(n8212), .A2(\srf/regTable[5][13] ), .B1(n8213), .B2(
        \srf/regTable[7][13] ), .ZN(n8269) );
  AOI22D1BWP U10575 ( .A1(n8210), .A2(\srf/regTable[4][13] ), .B1(n8211), .B2(
        \srf/regTable[6][13] ), .ZN(n8268) );
  AOI22D1BWP U10576 ( .A1(n8207), .A2(\srf/regTable[1][13] ), .B1(n8209), .B2(
        \srf/regTable[3][13] ), .ZN(n8267) );
  AOI22D1BWP U10577 ( .A1(n8203), .A2(\srf/regTable[0][13] ), .B1(n8205), .B2(
        \srf/regTable[2][13] ), .ZN(n8266) );
  ND4D1BWP U10578 ( .A1(n6136), .A2(n6137), .A3(n6138), .A4(n6139), .ZN(
        vectorData2[13]) );
  AOI22D1BWP U10579 ( .A1(n3569), .A2(\vrf/regTable[5][13] ), .B1(n3592), .B2(
        \vrf/regTable[7][13] ), .ZN(n6139) );
  AOI22D1BWP U10580 ( .A1(n3577), .A2(\vrf/regTable[4][13] ), .B1(n3591), .B2(
        \vrf/regTable[6][13] ), .ZN(n6138) );
  AOI22D1BWP U10581 ( .A1(n3571), .A2(\vrf/regTable[1][13] ), .B1(n3568), .B2(
        \vrf/regTable[3][13] ), .ZN(n6137) );
  AOI22D1BWP U10582 ( .A1(n3580), .A2(\vrf/regTable[0][13] ), .B1(n3566), .B2(
        \vrf/regTable[2][13] ), .ZN(n6136) );
  ND3D1BWP U10583 ( .A1(n5870), .A2(n5869), .A3(n5868), .ZN(n5871) );
  AOI211XD0BWP U10584 ( .A1(n5985), .A2(vectorData2[45]), .B(n5867), .C(n5866), 
        .ZN(n5868) );
  ND4D1BWP U10585 ( .A1(n5865), .A2(n5864), .A3(n5863), .A4(n5862), .ZN(n5866)
         );
  AOI22D1BWP U10586 ( .A1(n5978), .A2(vectorData2[205]), .B1(n5984), .B2(
        vectorData2[221]), .ZN(n5862) );
  ND4D1BWP U10587 ( .A1(n6968), .A2(n6969), .A3(n6970), .A4(n6971), .ZN(
        vectorData2[221]) );
  AOI22D1BWP U10588 ( .A1(n3569), .A2(\vrf/regTable[5][221] ), .B1(n3578), 
        .B2(\vrf/regTable[7][221] ), .ZN(n6971) );
  AOI22D1BWP U10589 ( .A1(n3577), .A2(\vrf/regTable[4][221] ), .B1(n3573), 
        .B2(\vrf/regTable[6][221] ), .ZN(n6970) );
  AOI22D1BWP U10590 ( .A1(n3571), .A2(\vrf/regTable[1][221] ), .B1(n3597), 
        .B2(\vrf/regTable[3][221] ), .ZN(n6969) );
  AOI22D1BWP U10591 ( .A1(n3580), .A2(\vrf/regTable[0][221] ), .B1(n3593), 
        .B2(\vrf/regTable[2][221] ), .ZN(n6968) );
  ND4D1BWP U10592 ( .A1(n6904), .A2(n6905), .A3(n6906), .A4(n6907), .ZN(
        vectorData2[205]) );
  AOI22D1BWP U10593 ( .A1(n3569), .A2(\vrf/regTable[5][205] ), .B1(n6083), 
        .B2(\vrf/regTable[7][205] ), .ZN(n6907) );
  AOI22D1BWP U10594 ( .A1(n3577), .A2(\vrf/regTable[4][205] ), .B1(n6081), 
        .B2(\vrf/regTable[6][205] ), .ZN(n6906) );
  AOI22D1BWP U10595 ( .A1(n3571), .A2(\vrf/regTable[1][205] ), .B1(n6079), 
        .B2(\vrf/regTable[3][205] ), .ZN(n6905) );
  AOI22D1BWP U10596 ( .A1(n3580), .A2(\vrf/regTable[0][205] ), .B1(n6075), 
        .B2(\vrf/regTable[2][205] ), .ZN(n6904) );
  AOI22D1BWP U10597 ( .A1(n5992), .A2(vectorData2[237]), .B1(n5976), .B2(
        vectorData2[109]), .ZN(n5863) );
  ND4D1BWP U10598 ( .A1(n6520), .A2(n6521), .A3(n6522), .A4(n6523), .ZN(
        vectorData2[109]) );
  AOI22D1BWP U10599 ( .A1(n3569), .A2(\vrf/regTable[5][109] ), .B1(n3578), 
        .B2(\vrf/regTable[7][109] ), .ZN(n6523) );
  AOI22D1BWP U10600 ( .A1(n8210), .A2(\vrf/regTable[4][109] ), .B1(n3573), 
        .B2(\vrf/regTable[6][109] ), .ZN(n6522) );
  AOI22D1BWP U10601 ( .A1(n3571), .A2(\vrf/regTable[1][109] ), .B1(n3597), 
        .B2(\vrf/regTable[3][109] ), .ZN(n6521) );
  AOI22D1BWP U10602 ( .A1(n8203), .A2(\vrf/regTable[0][109] ), .B1(n3593), 
        .B2(\vrf/regTable[2][109] ), .ZN(n6520) );
  ND4D1BWP U10603 ( .A1(n7032), .A2(n7033), .A3(n7034), .A4(n7035), .ZN(
        vectorData2[237]) );
  AOI22D1BWP U10604 ( .A1(n3569), .A2(\vrf/regTable[5][237] ), .B1(n3578), 
        .B2(\vrf/regTable[7][237] ), .ZN(n7035) );
  AOI22D1BWP U10605 ( .A1(n6080), .A2(\vrf/regTable[4][237] ), .B1(n3573), 
        .B2(\vrf/regTable[6][237] ), .ZN(n7034) );
  AOI22D1BWP U10606 ( .A1(n3571), .A2(\vrf/regTable[1][237] ), .B1(n3597), 
        .B2(\vrf/regTable[3][237] ), .ZN(n7033) );
  AOI22D1BWP U10607 ( .A1(n6073), .A2(\vrf/regTable[0][237] ), .B1(n3593), 
        .B2(\vrf/regTable[2][237] ), .ZN(n7032) );
  AOI22D1BWP U10608 ( .A1(n5974), .A2(vectorData2[61]), .B1(n5983), .B2(
        vectorData2[157]), .ZN(n5864) );
  ND4D1BWP U10609 ( .A1(n6712), .A2(n6713), .A3(n6714), .A4(n6715), .ZN(
        vectorData2[157]) );
  AOI22D1BWP U10610 ( .A1(n3569), .A2(\vrf/regTable[5][157] ), .B1(n3578), 
        .B2(\vrf/regTable[7][157] ), .ZN(n6715) );
  AOI22D1BWP U10611 ( .A1(n3577), .A2(\vrf/regTable[4][157] ), .B1(n3573), 
        .B2(\vrf/regTable[6][157] ), .ZN(n6714) );
  AOI22D1BWP U10612 ( .A1(n3571), .A2(\vrf/regTable[1][157] ), .B1(n3597), 
        .B2(\vrf/regTable[3][157] ), .ZN(n6713) );
  AOI22D1BWP U10613 ( .A1(n3580), .A2(\vrf/regTable[0][157] ), .B1(n3593), 
        .B2(\vrf/regTable[2][157] ), .ZN(n6712) );
  ND4D1BWP U10614 ( .A1(n6328), .A2(n6329), .A3(n6330), .A4(n6331), .ZN(
        vectorData2[61]) );
  AOI22D1BWP U10615 ( .A1(n3569), .A2(\vrf/regTable[5][61] ), .B1(n3592), .B2(
        \vrf/regTable[7][61] ), .ZN(n6331) );
  AOI22D1BWP U10616 ( .A1(n3577), .A2(\vrf/regTable[4][61] ), .B1(n3591), .B2(
        \vrf/regTable[6][61] ), .ZN(n6330) );
  AOI22D1BWP U10617 ( .A1(n3571), .A2(\vrf/regTable[1][61] ), .B1(n3568), .B2(
        \vrf/regTable[3][61] ), .ZN(n6329) );
  AOI22D1BWP U10618 ( .A1(n3580), .A2(\vrf/regTable[0][61] ), .B1(n3566), .B2(
        \vrf/regTable[2][61] ), .ZN(n6328) );
  AOI22D1BWP U10619 ( .A1(n5982), .A2(vectorData2[29]), .B1(n5980), .B2(
        vectorData2[253]), .ZN(n5865) );
  ND4D1BWP U10620 ( .A1(n7096), .A2(n7097), .A3(n7098), .A4(n7099), .ZN(
        vectorData2[253]) );
  AOI22D1BWP U10621 ( .A1(n3569), .A2(\vrf/regTable[5][253] ), .B1(n3578), 
        .B2(\vrf/regTable[7][253] ), .ZN(n7099) );
  AOI22D1BWP U10622 ( .A1(n3577), .A2(\vrf/regTable[4][253] ), .B1(n3573), 
        .B2(\vrf/regTable[6][253] ), .ZN(n7098) );
  AOI22D1BWP U10623 ( .A1(n3571), .A2(\vrf/regTable[1][253] ), .B1(n3597), 
        .B2(\vrf/regTable[3][253] ), .ZN(n7097) );
  AOI22D1BWP U10624 ( .A1(n3580), .A2(\vrf/regTable[0][253] ), .B1(n3593), 
        .B2(\vrf/regTable[2][253] ), .ZN(n7096) );
  ND4D1BWP U10625 ( .A1(n6200), .A2(n6201), .A3(n6202), .A4(n6203), .ZN(
        vectorData2[29]) );
  AOI22D1BWP U10626 ( .A1(n3569), .A2(\vrf/regTable[5][29] ), .B1(n3578), .B2(
        \vrf/regTable[7][29] ), .ZN(n6203) );
  AOI22D1BWP U10627 ( .A1(n3577), .A2(\vrf/regTable[4][29] ), .B1(n3573), .B2(
        \vrf/regTable[6][29] ), .ZN(n6202) );
  AOI22D1BWP U10628 ( .A1(n3571), .A2(\vrf/regTable[1][29] ), .B1(n3597), .B2(
        \vrf/regTable[3][29] ), .ZN(n6201) );
  AOI22D1BWP U10629 ( .A1(n3580), .A2(\vrf/regTable[0][29] ), .B1(n3593), .B2(
        \vrf/regTable[2][29] ), .ZN(n6200) );
  AO22D1BWP U10630 ( .A1(n5975), .A2(vectorData2[173]), .B1(n5977), .B2(
        vectorData2[141]), .Z(n5867) );
  ND4D1BWP U10631 ( .A1(n6648), .A2(n6649), .A3(n6650), .A4(n6651), .ZN(
        vectorData2[141]) );
  AOI22D1BWP U10632 ( .A1(n3569), .A2(\vrf/regTable[5][141] ), .B1(n3592), 
        .B2(\vrf/regTable[7][141] ), .ZN(n6651) );
  AOI22D1BWP U10633 ( .A1(n8210), .A2(\vrf/regTable[4][141] ), .B1(n3591), 
        .B2(\vrf/regTable[6][141] ), .ZN(n6650) );
  AOI22D1BWP U10634 ( .A1(n3571), .A2(\vrf/regTable[1][141] ), .B1(n3568), 
        .B2(\vrf/regTable[3][141] ), .ZN(n6649) );
  AOI22D1BWP U10635 ( .A1(n8203), .A2(\vrf/regTable[0][141] ), .B1(n3566), 
        .B2(\vrf/regTable[2][141] ), .ZN(n6648) );
  ND4D1BWP U10636 ( .A1(n6776), .A2(n6777), .A3(n6778), .A4(n6779), .ZN(
        vectorData2[173]) );
  AOI22D1BWP U10637 ( .A1(n3569), .A2(\vrf/regTable[5][173] ), .B1(n6083), 
        .B2(\vrf/regTable[7][173] ), .ZN(n6779) );
  AOI22D1BWP U10638 ( .A1(n3577), .A2(\vrf/regTable[4][173] ), .B1(n6081), 
        .B2(\vrf/regTable[6][173] ), .ZN(n6778) );
  AOI22D1BWP U10639 ( .A1(n3571), .A2(\vrf/regTable[1][173] ), .B1(n6079), 
        .B2(\vrf/regTable[3][173] ), .ZN(n6777) );
  AOI22D1BWP U10640 ( .A1(n3580), .A2(\vrf/regTable[0][173] ), .B1(n6075), 
        .B2(\vrf/regTable[2][173] ), .ZN(n6776) );
  ND4D1BWP U10641 ( .A1(n6264), .A2(n6265), .A3(n6266), .A4(n6267), .ZN(
        vectorData2[45]) );
  AOI22D1BWP U10642 ( .A1(n3569), .A2(\vrf/regTable[5][45] ), .B1(n3578), .B2(
        \vrf/regTable[7][45] ), .ZN(n6267) );
  AOI22D1BWP U10643 ( .A1(n3577), .A2(\vrf/regTable[4][45] ), .B1(n3573), .B2(
        \vrf/regTable[6][45] ), .ZN(n6266) );
  AOI22D1BWP U10644 ( .A1(n3571), .A2(\vrf/regTable[1][45] ), .B1(n3597), .B2(
        \vrf/regTable[3][45] ), .ZN(n6265) );
  AOI22D1BWP U10645 ( .A1(n3580), .A2(\vrf/regTable[0][45] ), .B1(n3593), .B2(
        \vrf/regTable[2][45] ), .ZN(n6264) );
  AOI22D1BWP U10646 ( .A1(n5981), .A2(vectorData2[189]), .B1(n5972), .B2(
        vectorData2[125]), .ZN(n5869) );
  ND4D1BWP U10647 ( .A1(n6584), .A2(n6585), .A3(n6586), .A4(n6587), .ZN(
        vectorData2[125]) );
  AOI22D1BWP U10648 ( .A1(n3569), .A2(\vrf/regTable[5][125] ), .B1(n3592), 
        .B2(\vrf/regTable[7][125] ), .ZN(n6587) );
  AOI22D1BWP U10649 ( .A1(n3577), .A2(\vrf/regTable[4][125] ), .B1(n3591), 
        .B2(\vrf/regTable[6][125] ), .ZN(n6586) );
  AOI22D1BWP U10650 ( .A1(n3571), .A2(\vrf/regTable[1][125] ), .B1(n3568), 
        .B2(\vrf/regTable[3][125] ), .ZN(n6585) );
  AOI22D1BWP U10651 ( .A1(n3580), .A2(\vrf/regTable[0][125] ), .B1(n3566), 
        .B2(\vrf/regTable[2][125] ), .ZN(n6584) );
  ND4D1BWP U10652 ( .A1(n6840), .A2(n6841), .A3(n6842), .A4(n6843), .ZN(
        vectorData2[189]) );
  AOI22D1BWP U10653 ( .A1(n3569), .A2(\vrf/regTable[5][189] ), .B1(n3592), 
        .B2(\vrf/regTable[7][189] ), .ZN(n6843) );
  AOI22D1BWP U10654 ( .A1(n3577), .A2(\vrf/regTable[4][189] ), .B1(n3591), 
        .B2(\vrf/regTable[6][189] ), .ZN(n6842) );
  AOI22D1BWP U10655 ( .A1(n3571), .A2(\vrf/regTable[1][189] ), .B1(n3568), 
        .B2(\vrf/regTable[3][189] ), .ZN(n6841) );
  AOI22D1BWP U10656 ( .A1(n3580), .A2(\vrf/regTable[0][189] ), .B1(n3566), 
        .B2(\vrf/regTable[2][189] ), .ZN(n6840) );
  AOI22D1BWP U10657 ( .A1(n5979), .A2(vectorData2[93]), .B1(n5973), .B2(
        vectorData2[77]), .ZN(n5870) );
  ND4D1BWP U10658 ( .A1(n6392), .A2(n6393), .A3(n6394), .A4(n6395), .ZN(
        vectorData2[77]) );
  AOI22D1BWP U10659 ( .A1(n3569), .A2(\vrf/regTable[5][77] ), .B1(n3578), .B2(
        \vrf/regTable[7][77] ), .ZN(n6395) );
  AOI22D1BWP U10660 ( .A1(n3577), .A2(\vrf/regTable[4][77] ), .B1(n3573), .B2(
        \vrf/regTable[6][77] ), .ZN(n6394) );
  AOI22D1BWP U10661 ( .A1(n3571), .A2(\vrf/regTable[1][77] ), .B1(n3597), .B2(
        \vrf/regTable[3][77] ), .ZN(n6393) );
  AOI22D1BWP U10662 ( .A1(n3580), .A2(\vrf/regTable[0][77] ), .B1(n3593), .B2(
        \vrf/regTable[2][77] ), .ZN(n6392) );
  ND4D1BWP U10663 ( .A1(n6456), .A2(n6457), .A3(n6458), .A4(n6459), .ZN(
        vectorData2[93]) );
  AOI22D1BWP U10664 ( .A1(n3569), .A2(\vrf/regTable[5][93] ), .B1(n3592), .B2(
        \vrf/regTable[7][93] ), .ZN(n6459) );
  AOI22D1BWP U10665 ( .A1(n3577), .A2(\vrf/regTable[4][93] ), .B1(n3591), .B2(
        \vrf/regTable[6][93] ), .ZN(n6458) );
  AOI22D1BWP U10666 ( .A1(n3571), .A2(\vrf/regTable[1][93] ), .B1(n3568), .B2(
        \vrf/regTable[3][93] ), .ZN(n6457) );
  AOI22D1BWP U10667 ( .A1(n3580), .A2(\vrf/regTable[0][93] ), .B1(n3566), .B2(
        \vrf/regTable[2][93] ), .ZN(n6456) );
  AO222D1BWP U10668 ( .A1(vectorData2[14]), .A2(n4570), .B1(n4569), .B2(
        scalarData2[14]), .C1(WR), .C2(n5881), .Z(dataOut[14]) );
  ND3D1BWP U10669 ( .A1(n5880), .A2(n5879), .A3(n5878), .ZN(n5881) );
  AOI211XD0BWP U10670 ( .A1(n5974), .A2(vectorData2[62]), .B(n5877), .C(n5876), 
        .ZN(n5878) );
  ND4D1BWP U10671 ( .A1(n5875), .A2(n5874), .A3(n5873), .A4(n5872), .ZN(n5876)
         );
  AOI22D1BWP U10672 ( .A1(n5980), .A2(vectorData2[254]), .B1(n5976), .B2(
        vectorData2[110]), .ZN(n5872) );
  ND4D1BWP U10673 ( .A1(n6524), .A2(n6525), .A3(n6526), .A4(n6527), .ZN(
        vectorData2[110]) );
  AOI22D1BWP U10674 ( .A1(n3569), .A2(\vrf/regTable[5][110] ), .B1(n3578), 
        .B2(\vrf/regTable[7][110] ), .ZN(n6527) );
  AOI22D1BWP U10675 ( .A1(n3577), .A2(\vrf/regTable[4][110] ), .B1(n3573), 
        .B2(\vrf/regTable[6][110] ), .ZN(n6526) );
  AOI22D1BWP U10676 ( .A1(n3571), .A2(\vrf/regTable[1][110] ), .B1(n3597), 
        .B2(\vrf/regTable[3][110] ), .ZN(n6525) );
  AOI22D1BWP U10677 ( .A1(n3580), .A2(\vrf/regTable[0][110] ), .B1(n3593), 
        .B2(\vrf/regTable[2][110] ), .ZN(n6524) );
  ND4D1BWP U10678 ( .A1(n7100), .A2(n7101), .A3(n7102), .A4(n7103), .ZN(
        vectorData2[254]) );
  AOI22D1BWP U10679 ( .A1(n3569), .A2(\vrf/regTable[5][254] ), .B1(n6083), 
        .B2(\vrf/regTable[7][254] ), .ZN(n7103) );
  AOI22D1BWP U10680 ( .A1(n3577), .A2(\vrf/regTable[4][254] ), .B1(n6081), 
        .B2(\vrf/regTable[6][254] ), .ZN(n7102) );
  AOI22D1BWP U10681 ( .A1(n3571), .A2(\vrf/regTable[1][254] ), .B1(n6079), 
        .B2(\vrf/regTable[3][254] ), .ZN(n7101) );
  AOI22D1BWP U10682 ( .A1(n3580), .A2(\vrf/regTable[0][254] ), .B1(n6075), 
        .B2(\vrf/regTable[2][254] ), .ZN(n7100) );
  AOI22D1BWP U10683 ( .A1(n5979), .A2(vectorData2[94]), .B1(n5992), .B2(
        vectorData2[238]), .ZN(n5873) );
  ND4D1BWP U10684 ( .A1(n7036), .A2(n7037), .A3(n7038), .A4(n7039), .ZN(
        vectorData2[238]) );
  AOI22D1BWP U10685 ( .A1(n3569), .A2(\vrf/regTable[5][238] ), .B1(n3578), 
        .B2(\vrf/regTable[7][238] ), .ZN(n7039) );
  AOI22D1BWP U10686 ( .A1(n3577), .A2(\vrf/regTable[4][238] ), .B1(n3573), 
        .B2(\vrf/regTable[6][238] ), .ZN(n7038) );
  AOI22D1BWP U10687 ( .A1(n3571), .A2(\vrf/regTable[1][238] ), .B1(n3597), 
        .B2(\vrf/regTable[3][238] ), .ZN(n7037) );
  AOI22D1BWP U10688 ( .A1(n3580), .A2(\vrf/regTable[0][238] ), .B1(n3593), 
        .B2(\vrf/regTable[2][238] ), .ZN(n7036) );
  ND4D1BWP U10689 ( .A1(n6460), .A2(n6461), .A3(n6462), .A4(n6463), .ZN(
        vectorData2[94]) );
  AOI22D1BWP U10690 ( .A1(n6082), .A2(\vrf/regTable[5][94] ), .B1(n3592), .B2(
        \vrf/regTable[7][94] ), .ZN(n6463) );
  AOI22D1BWP U10691 ( .A1(n6080), .A2(\vrf/regTable[4][94] ), .B1(n3591), .B2(
        \vrf/regTable[6][94] ), .ZN(n6462) );
  AOI22D1BWP U10692 ( .A1(n6077), .A2(\vrf/regTable[1][94] ), .B1(n3568), .B2(
        \vrf/regTable[3][94] ), .ZN(n6461) );
  AOI22D1BWP U10693 ( .A1(n6073), .A2(\vrf/regTable[0][94] ), .B1(n3566), .B2(
        \vrf/regTable[2][94] ), .ZN(n6460) );
  AOI22D1BWP U10694 ( .A1(n5975), .A2(vectorData2[174]), .B1(n5983), .B2(
        vectorData2[158]), .ZN(n5874) );
  ND4D1BWP U10695 ( .A1(n6716), .A2(n6717), .A3(n6718), .A4(n6719), .ZN(
        vectorData2[158]) );
  AOI22D1BWP U10696 ( .A1(n3569), .A2(\vrf/regTable[5][158] ), .B1(n3592), 
        .B2(\vrf/regTable[7][158] ), .ZN(n6719) );
  AOI22D1BWP U10697 ( .A1(n3577), .A2(\vrf/regTable[4][158] ), .B1(n3591), 
        .B2(\vrf/regTable[6][158] ), .ZN(n6718) );
  AOI22D1BWP U10698 ( .A1(n3571), .A2(\vrf/regTable[1][158] ), .B1(n3568), 
        .B2(\vrf/regTable[3][158] ), .ZN(n6717) );
  AOI22D1BWP U10699 ( .A1(n3580), .A2(\vrf/regTable[0][158] ), .B1(n3566), 
        .B2(\vrf/regTable[2][158] ), .ZN(n6716) );
  ND4D1BWP U10700 ( .A1(n6780), .A2(n6781), .A3(n6782), .A4(n6783), .ZN(
        vectorData2[174]) );
  AOI22D1BWP U10701 ( .A1(n3569), .A2(\vrf/regTable[5][174] ), .B1(n3578), 
        .B2(\vrf/regTable[7][174] ), .ZN(n6783) );
  AOI22D1BWP U10702 ( .A1(n3577), .A2(\vrf/regTable[4][174] ), .B1(n3573), 
        .B2(\vrf/regTable[6][174] ), .ZN(n6782) );
  AOI22D1BWP U10703 ( .A1(n3571), .A2(\vrf/regTable[1][174] ), .B1(n3597), 
        .B2(\vrf/regTable[3][174] ), .ZN(n6781) );
  AOI22D1BWP U10704 ( .A1(n3580), .A2(\vrf/regTable[0][174] ), .B1(n3593), 
        .B2(\vrf/regTable[2][174] ), .ZN(n6780) );
  AOI22D1BWP U10705 ( .A1(n5981), .A2(vectorData2[190]), .B1(n5978), .B2(
        vectorData2[206]), .ZN(n5875) );
  ND4D1BWP U10706 ( .A1(n6908), .A2(n6909), .A3(n6910), .A4(n6911), .ZN(
        vectorData2[206]) );
  AOI22D1BWP U10707 ( .A1(n3569), .A2(\vrf/regTable[5][206] ), .B1(n3592), 
        .B2(\vrf/regTable[7][206] ), .ZN(n6911) );
  AOI22D1BWP U10708 ( .A1(n3577), .A2(\vrf/regTable[4][206] ), .B1(n3591), 
        .B2(\vrf/regTable[6][206] ), .ZN(n6910) );
  AOI22D1BWP U10709 ( .A1(n3571), .A2(\vrf/regTable[1][206] ), .B1(n3568), 
        .B2(\vrf/regTable[3][206] ), .ZN(n6909) );
  AOI22D1BWP U10710 ( .A1(n3580), .A2(\vrf/regTable[0][206] ), .B1(n3566), 
        .B2(\vrf/regTable[2][206] ), .ZN(n6908) );
  ND4D1BWP U10711 ( .A1(n6844), .A2(n6845), .A3(n6846), .A4(n6847), .ZN(
        vectorData2[190]) );
  AOI22D1BWP U10712 ( .A1(n3569), .A2(\vrf/regTable[5][190] ), .B1(n3578), 
        .B2(\vrf/regTable[7][190] ), .ZN(n6847) );
  AOI22D1BWP U10713 ( .A1(n3577), .A2(\vrf/regTable[4][190] ), .B1(n3573), 
        .B2(\vrf/regTable[6][190] ), .ZN(n6846) );
  AOI22D1BWP U10714 ( .A1(n3571), .A2(\vrf/regTable[1][190] ), .B1(n3597), 
        .B2(\vrf/regTable[3][190] ), .ZN(n6845) );
  AOI22D1BWP U10715 ( .A1(n3580), .A2(\vrf/regTable[0][190] ), .B1(n3593), 
        .B2(\vrf/regTable[2][190] ), .ZN(n6844) );
  AO22D1BWP U10716 ( .A1(n5973), .A2(vectorData2[78]), .B1(n5972), .B2(
        vectorData2[126]), .Z(n5877) );
  ND4D1BWP U10717 ( .A1(n6588), .A2(n6589), .A3(n6590), .A4(n6591), .ZN(
        vectorData2[126]) );
  AOI22D1BWP U10718 ( .A1(n3569), .A2(\vrf/regTable[5][126] ), .B1(n3592), 
        .B2(\vrf/regTable[7][126] ), .ZN(n6591) );
  AOI22D1BWP U10719 ( .A1(n3577), .A2(\vrf/regTable[4][126] ), .B1(n3591), 
        .B2(\vrf/regTable[6][126] ), .ZN(n6590) );
  AOI22D1BWP U10720 ( .A1(n3571), .A2(\vrf/regTable[1][126] ), .B1(n3568), 
        .B2(\vrf/regTable[3][126] ), .ZN(n6589) );
  AOI22D1BWP U10721 ( .A1(n3580), .A2(\vrf/regTable[0][126] ), .B1(n3566), 
        .B2(\vrf/regTable[2][126] ), .ZN(n6588) );
  ND4D1BWP U10722 ( .A1(n6396), .A2(n6397), .A3(n6398), .A4(n6399), .ZN(
        vectorData2[78]) );
  AOI22D1BWP U10723 ( .A1(n6082), .A2(\vrf/regTable[5][78] ), .B1(n3578), .B2(
        \vrf/regTable[7][78] ), .ZN(n6399) );
  AOI22D1BWP U10724 ( .A1(n6080), .A2(\vrf/regTable[4][78] ), .B1(n3573), .B2(
        \vrf/regTable[6][78] ), .ZN(n6398) );
  AOI22D1BWP U10725 ( .A1(n6077), .A2(\vrf/regTable[1][78] ), .B1(n3597), .B2(
        \vrf/regTable[3][78] ), .ZN(n6397) );
  AOI22D1BWP U10726 ( .A1(n6073), .A2(\vrf/regTable[0][78] ), .B1(n3593), .B2(
        \vrf/regTable[2][78] ), .ZN(n6396) );
  ND4D1BWP U10727 ( .A1(n6332), .A2(n6333), .A3(n6334), .A4(n6335), .ZN(
        vectorData2[62]) );
  AOI22D1BWP U10728 ( .A1(n3569), .A2(\vrf/regTable[5][62] ), .B1(n3592), .B2(
        \vrf/regTable[7][62] ), .ZN(n6335) );
  AOI22D1BWP U10729 ( .A1(n3577), .A2(\vrf/regTable[4][62] ), .B1(n3591), .B2(
        \vrf/regTable[6][62] ), .ZN(n6334) );
  AOI22D1BWP U10730 ( .A1(n3571), .A2(\vrf/regTable[1][62] ), .B1(n3568), .B2(
        \vrf/regTable[3][62] ), .ZN(n6333) );
  AOI22D1BWP U10731 ( .A1(n3580), .A2(\vrf/regTable[0][62] ), .B1(n3566), .B2(
        \vrf/regTable[2][62] ), .ZN(n6332) );
  AOI22D1BWP U10732 ( .A1(n5977), .A2(vectorData2[142]), .B1(n5982), .B2(
        vectorData2[30]), .ZN(n5879) );
  ND4D1BWP U10733 ( .A1(n6204), .A2(n6205), .A3(n6206), .A4(n6207), .ZN(
        vectorData2[30]) );
  AOI22D1BWP U10734 ( .A1(n3569), .A2(\vrf/regTable[5][30] ), .B1(n3592), .B2(
        \vrf/regTable[7][30] ), .ZN(n6207) );
  AOI22D1BWP U10735 ( .A1(n3577), .A2(\vrf/regTable[4][30] ), .B1(n3591), .B2(
        \vrf/regTable[6][30] ), .ZN(n6206) );
  AOI22D1BWP U10736 ( .A1(n3571), .A2(\vrf/regTable[1][30] ), .B1(n3568), .B2(
        \vrf/regTable[3][30] ), .ZN(n6205) );
  AOI22D1BWP U10737 ( .A1(n3580), .A2(\vrf/regTable[0][30] ), .B1(n3566), .B2(
        \vrf/regTable[2][30] ), .ZN(n6204) );
  ND4D1BWP U10738 ( .A1(n6652), .A2(n6653), .A3(n6654), .A4(n6655), .ZN(
        vectorData2[142]) );
  AOI22D1BWP U10739 ( .A1(n3569), .A2(\vrf/regTable[5][142] ), .B1(n3578), 
        .B2(\vrf/regTable[7][142] ), .ZN(n6655) );
  AOI22D1BWP U10740 ( .A1(n3577), .A2(\vrf/regTable[4][142] ), .B1(n3573), 
        .B2(\vrf/regTable[6][142] ), .ZN(n6654) );
  AOI22D1BWP U10741 ( .A1(n3571), .A2(\vrf/regTable[1][142] ), .B1(n3597), 
        .B2(\vrf/regTable[3][142] ), .ZN(n6653) );
  AOI22D1BWP U10742 ( .A1(n3580), .A2(\vrf/regTable[0][142] ), .B1(n3593), 
        .B2(\vrf/regTable[2][142] ), .ZN(n6652) );
  AOI22D1BWP U10743 ( .A1(n5985), .A2(vectorData2[46]), .B1(n5984), .B2(
        vectorData2[222]), .ZN(n5880) );
  ND4D1BWP U10744 ( .A1(n6972), .A2(n6973), .A3(n6974), .A4(n6975), .ZN(
        vectorData2[222]) );
  AOI22D1BWP U10745 ( .A1(n3569), .A2(\vrf/regTable[5][222] ), .B1(n3578), 
        .B2(\vrf/regTable[7][222] ), .ZN(n6975) );
  AOI22D1BWP U10746 ( .A1(n3577), .A2(\vrf/regTable[4][222] ), .B1(n3573), 
        .B2(\vrf/regTable[6][222] ), .ZN(n6974) );
  AOI22D1BWP U10747 ( .A1(n3571), .A2(\vrf/regTable[1][222] ), .B1(n3597), 
        .B2(\vrf/regTable[3][222] ), .ZN(n6973) );
  AOI22D1BWP U10748 ( .A1(n3580), .A2(\vrf/regTable[0][222] ), .B1(n3593), 
        .B2(\vrf/regTable[2][222] ), .ZN(n6972) );
  ND4D1BWP U10749 ( .A1(n6268), .A2(n6269), .A3(n6270), .A4(n6271), .ZN(
        vectorData2[46]) );
  AOI22D1BWP U10750 ( .A1(n3569), .A2(\vrf/regTable[5][46] ), .B1(n3578), .B2(
        \vrf/regTable[7][46] ), .ZN(n6271) );
  AOI22D1BWP U10751 ( .A1(n3577), .A2(\vrf/regTable[4][46] ), .B1(n3573), .B2(
        \vrf/regTable[6][46] ), .ZN(n6270) );
  AOI22D1BWP U10752 ( .A1(n3571), .A2(\vrf/regTable[1][46] ), .B1(n3597), .B2(
        \vrf/regTable[3][46] ), .ZN(n6269) );
  AOI22D1BWP U10753 ( .A1(n3580), .A2(\vrf/regTable[0][46] ), .B1(n3593), .B2(
        \vrf/regTable[2][46] ), .ZN(n6268) );
  ND4D1BWP U10754 ( .A1(n8270), .A2(n8271), .A3(n8272), .A4(n8273), .ZN(
        scalarData2[14]) );
  AOI22D1BWP U10755 ( .A1(n8212), .A2(\srf/regTable[5][14] ), .B1(n8213), .B2(
        \srf/regTable[7][14] ), .ZN(n8273) );
  AOI22D1BWP U10756 ( .A1(n8210), .A2(\srf/regTable[4][14] ), .B1(n8211), .B2(
        \srf/regTable[6][14] ), .ZN(n8272) );
  AOI22D1BWP U10757 ( .A1(n8207), .A2(\srf/regTable[1][14] ), .B1(n8209), .B2(
        \srf/regTable[3][14] ), .ZN(n8271) );
  AOI22D1BWP U10758 ( .A1(n8203), .A2(\srf/regTable[0][14] ), .B1(n8205), .B2(
        \srf/regTable[2][14] ), .ZN(n8270) );
  ND4D1BWP U10759 ( .A1(n6140), .A2(n6141), .A3(n6142), .A4(n6143), .ZN(
        vectorData2[14]) );
  AOI22D1BWP U10760 ( .A1(n3569), .A2(\vrf/regTable[5][14] ), .B1(n3592), .B2(
        \vrf/regTable[7][14] ), .ZN(n6143) );
  AOI22D1BWP U10761 ( .A1(n3577), .A2(\vrf/regTable[4][14] ), .B1(n3591), .B2(
        \vrf/regTable[6][14] ), .ZN(n6142) );
  AOI22D1BWP U10762 ( .A1(n3571), .A2(\vrf/regTable[1][14] ), .B1(n3568), .B2(
        \vrf/regTable[3][14] ), .ZN(n6141) );
  AOI22D1BWP U10763 ( .A1(n3580), .A2(\vrf/regTable[0][14] ), .B1(n3566), .B2(
        \vrf/regTable[2][14] ), .ZN(n6140) );
  AO222D1BWP U10764 ( .A1(WR), .A2(n5891), .B1(n4570), .B2(vectorData2[15]), 
        .C1(n4569), .C2(scalarData2[15]), .Z(dataOut[15]) );
  ND4D1BWP U10765 ( .A1(n8274), .A2(n8275), .A3(n8276), .A4(n8277), .ZN(
        scalarData2[15]) );
  AOI22D1BWP U10766 ( .A1(n8212), .A2(\srf/regTable[5][15] ), .B1(n8213), .B2(
        \srf/regTable[7][15] ), .ZN(n8277) );
  AOI22D1BWP U10767 ( .A1(n8210), .A2(\srf/regTable[4][15] ), .B1(n8211), .B2(
        \srf/regTable[6][15] ), .ZN(n8276) );
  AOI22D1BWP U10768 ( .A1(n8207), .A2(\srf/regTable[1][15] ), .B1(n8209), .B2(
        \srf/regTable[3][15] ), .ZN(n8275) );
  AOI22D1BWP U10769 ( .A1(n8203), .A2(\srf/regTable[0][15] ), .B1(n8205), .B2(
        \srf/regTable[2][15] ), .ZN(n8274) );
  ND4D1BWP U10770 ( .A1(n6144), .A2(n6145), .A3(n6146), .A4(n6147), .ZN(
        vectorData2[15]) );
  AOI22D1BWP U10771 ( .A1(n3569), .A2(\vrf/regTable[5][15] ), .B1(n3592), .B2(
        \vrf/regTable[7][15] ), .ZN(n6147) );
  AOI22D1BWP U10772 ( .A1(n3577), .A2(\vrf/regTable[4][15] ), .B1(n3591), .B2(
        \vrf/regTable[6][15] ), .ZN(n6146) );
  AOI22D1BWP U10773 ( .A1(n3571), .A2(\vrf/regTable[1][15] ), .B1(n3568), .B2(
        \vrf/regTable[3][15] ), .ZN(n6145) );
  AOI22D1BWP U10774 ( .A1(n3580), .A2(\vrf/regTable[0][15] ), .B1(n3566), .B2(
        \vrf/regTable[2][15] ), .ZN(n6144) );
  ND3D1BWP U10775 ( .A1(n5890), .A2(n5889), .A3(n5888), .ZN(n5891) );
  AOI211XD0BWP U10776 ( .A1(n5981), .A2(vectorData2[191]), .B(n5887), .C(n5886), .ZN(n5888) );
  ND4D1BWP U10777 ( .A1(n5885), .A2(n5884), .A3(n5883), .A4(n5882), .ZN(n5886)
         );
  AOI22D1BWP U10778 ( .A1(n5978), .A2(vectorData2[207]), .B1(n5980), .B2(
        vectorData2[255]), .ZN(n5882) );
  ND4D1BWP U10779 ( .A1(n7104), .A2(n7105), .A3(n7106), .A4(n7107), .ZN(
        vectorData2[255]) );
  AOI22D1BWP U10780 ( .A1(n3569), .A2(\vrf/regTable[5][255] ), .B1(n3592), 
        .B2(\vrf/regTable[7][255] ), .ZN(n7107) );
  AOI22D1BWP U10781 ( .A1(n3577), .A2(\vrf/regTable[4][255] ), .B1(n3591), 
        .B2(\vrf/regTable[6][255] ), .ZN(n7106) );
  AOI22D1BWP U10782 ( .A1(n3571), .A2(\vrf/regTable[1][255] ), .B1(n3568), 
        .B2(\vrf/regTable[3][255] ), .ZN(n7105) );
  AOI22D1BWP U10783 ( .A1(n3580), .A2(\vrf/regTable[0][255] ), .B1(n3566), 
        .B2(\vrf/regTable[2][255] ), .ZN(n7104) );
  ND4D1BWP U10784 ( .A1(n6912), .A2(n6913), .A3(n6914), .A4(n6915), .ZN(
        vectorData2[207]) );
  AOI22D1BWP U10785 ( .A1(n3569), .A2(\vrf/regTable[5][207] ), .B1(n3578), 
        .B2(\vrf/regTable[7][207] ), .ZN(n6915) );
  AOI22D1BWP U10786 ( .A1(n3577), .A2(\vrf/regTable[4][207] ), .B1(n3573), 
        .B2(\vrf/regTable[6][207] ), .ZN(n6914) );
  AOI22D1BWP U10787 ( .A1(n3571), .A2(\vrf/regTable[1][207] ), .B1(n3597), 
        .B2(\vrf/regTable[3][207] ), .ZN(n6913) );
  AOI22D1BWP U10788 ( .A1(n3580), .A2(\vrf/regTable[0][207] ), .B1(n3593), 
        .B2(\vrf/regTable[2][207] ), .ZN(n6912) );
  AOI22D1BWP U10789 ( .A1(n5985), .A2(vectorData2[47]), .B1(n5976), .B2(
        vectorData2[111]), .ZN(n5883) );
  ND4D1BWP U10790 ( .A1(n6528), .A2(n6529), .A3(n6530), .A4(n6531), .ZN(
        vectorData2[111]) );
  AOI22D1BWP U10791 ( .A1(n3569), .A2(\vrf/regTable[5][111] ), .B1(n3578), 
        .B2(\vrf/regTable[7][111] ), .ZN(n6531) );
  AOI22D1BWP U10792 ( .A1(n6080), .A2(\vrf/regTable[4][111] ), .B1(n3573), 
        .B2(\vrf/regTable[6][111] ), .ZN(n6530) );
  AOI22D1BWP U10793 ( .A1(n3571), .A2(\vrf/regTable[1][111] ), .B1(n3597), 
        .B2(\vrf/regTable[3][111] ), .ZN(n6529) );
  AOI22D1BWP U10794 ( .A1(n6073), .A2(\vrf/regTable[0][111] ), .B1(n3593), 
        .B2(\vrf/regTable[2][111] ), .ZN(n6528) );
  ND4D1BWP U10795 ( .A1(n6272), .A2(n6273), .A3(n6274), .A4(n6275), .ZN(
        vectorData2[47]) );
  AOI22D1BWP U10796 ( .A1(n3569), .A2(\vrf/regTable[5][47] ), .B1(n3578), .B2(
        \vrf/regTable[7][47] ), .ZN(n6275) );
  AOI22D1BWP U10797 ( .A1(n3577), .A2(\vrf/regTable[4][47] ), .B1(n3573), .B2(
        \vrf/regTable[6][47] ), .ZN(n6274) );
  AOI22D1BWP U10798 ( .A1(n3571), .A2(\vrf/regTable[1][47] ), .B1(n3597), .B2(
        \vrf/regTable[3][47] ), .ZN(n6273) );
  AOI22D1BWP U10799 ( .A1(n3580), .A2(\vrf/regTable[0][47] ), .B1(n3593), .B2(
        \vrf/regTable[2][47] ), .ZN(n6272) );
  AOI22D1BWP U10800 ( .A1(n5979), .A2(vectorData2[95]), .B1(n5992), .B2(
        vectorData2[239]), .ZN(n5884) );
  ND4D1BWP U10801 ( .A1(n7040), .A2(n7041), .A3(n7042), .A4(n7043), .ZN(
        vectorData2[239]) );
  AOI22D1BWP U10802 ( .A1(n3569), .A2(\vrf/regTable[5][239] ), .B1(n3578), 
        .B2(\vrf/regTable[7][239] ), .ZN(n7043) );
  AOI22D1BWP U10803 ( .A1(n3577), .A2(\vrf/regTable[4][239] ), .B1(n3573), 
        .B2(\vrf/regTable[6][239] ), .ZN(n7042) );
  AOI22D1BWP U10804 ( .A1(n3571), .A2(\vrf/regTable[1][239] ), .B1(n3597), 
        .B2(\vrf/regTable[3][239] ), .ZN(n7041) );
  AOI22D1BWP U10805 ( .A1(n3580), .A2(\vrf/regTable[0][239] ), .B1(n3593), 
        .B2(\vrf/regTable[2][239] ), .ZN(n7040) );
  ND4D1BWP U10806 ( .A1(n6464), .A2(n6465), .A3(n6466), .A4(n6467), .ZN(
        vectorData2[95]) );
  AOI22D1BWP U10807 ( .A1(n3569), .A2(\vrf/regTable[5][95] ), .B1(n3592), .B2(
        \vrf/regTable[7][95] ), .ZN(n6467) );
  AOI22D1BWP U10808 ( .A1(n3577), .A2(\vrf/regTable[4][95] ), .B1(n3591), .B2(
        \vrf/regTable[6][95] ), .ZN(n6466) );
  AOI22D1BWP U10809 ( .A1(n3571), .A2(\vrf/regTable[1][95] ), .B1(n3568), .B2(
        \vrf/regTable[3][95] ), .ZN(n6465) );
  AOI22D1BWP U10810 ( .A1(n3580), .A2(\vrf/regTable[0][95] ), .B1(n3566), .B2(
        \vrf/regTable[2][95] ), .ZN(n6464) );
  AOI22D1BWP U10811 ( .A1(n5973), .A2(vectorData2[79]), .B1(n5983), .B2(
        vectorData2[159]), .ZN(n5885) );
  ND4D1BWP U10812 ( .A1(n6720), .A2(n6721), .A3(n6722), .A4(n6723), .ZN(
        vectorData2[159]) );
  AOI22D1BWP U10813 ( .A1(n3569), .A2(\vrf/regTable[5][159] ), .B1(n3578), 
        .B2(\vrf/regTable[7][159] ), .ZN(n6723) );
  AOI22D1BWP U10814 ( .A1(n3577), .A2(\vrf/regTable[4][159] ), .B1(n3573), 
        .B2(\vrf/regTable[6][159] ), .ZN(n6722) );
  AOI22D1BWP U10815 ( .A1(n3571), .A2(\vrf/regTable[1][159] ), .B1(n3597), 
        .B2(\vrf/regTable[3][159] ), .ZN(n6721) );
  AOI22D1BWP U10816 ( .A1(n3580), .A2(\vrf/regTable[0][159] ), .B1(n3593), 
        .B2(\vrf/regTable[2][159] ), .ZN(n6720) );
  ND4D1BWP U10817 ( .A1(n6400), .A2(n6401), .A3(n6402), .A4(n6403), .ZN(
        vectorData2[79]) );
  AOI22D1BWP U10818 ( .A1(n3569), .A2(\vrf/regTable[5][79] ), .B1(n3592), .B2(
        \vrf/regTable[7][79] ), .ZN(n6403) );
  AOI22D1BWP U10819 ( .A1(n3577), .A2(\vrf/regTable[4][79] ), .B1(n3591), .B2(
        \vrf/regTable[6][79] ), .ZN(n6402) );
  AOI22D1BWP U10820 ( .A1(n3571), .A2(\vrf/regTable[1][79] ), .B1(n3568), .B2(
        \vrf/regTable[3][79] ), .ZN(n6401) );
  AOI22D1BWP U10821 ( .A1(n3580), .A2(\vrf/regTable[0][79] ), .B1(n3566), .B2(
        \vrf/regTable[2][79] ), .ZN(n6400) );
  AO22D1BWP U10822 ( .A1(n5974), .A2(vectorData2[63]), .B1(n5972), .B2(
        vectorData2[127]), .Z(n5887) );
  ND4D1BWP U10823 ( .A1(n6592), .A2(n6593), .A3(n6594), .A4(n6595), .ZN(
        vectorData2[127]) );
  AOI22D1BWP U10824 ( .A1(n3569), .A2(\vrf/regTable[5][127] ), .B1(n3592), 
        .B2(\vrf/regTable[7][127] ), .ZN(n6595) );
  AOI22D1BWP U10825 ( .A1(n3577), .A2(\vrf/regTable[4][127] ), .B1(n3591), 
        .B2(\vrf/regTable[6][127] ), .ZN(n6594) );
  AOI22D1BWP U10826 ( .A1(n3571), .A2(\vrf/regTable[1][127] ), .B1(n3568), 
        .B2(\vrf/regTable[3][127] ), .ZN(n6593) );
  AOI22D1BWP U10827 ( .A1(n3580), .A2(\vrf/regTable[0][127] ), .B1(n3566), 
        .B2(\vrf/regTable[2][127] ), .ZN(n6592) );
  ND4D1BWP U10828 ( .A1(n6336), .A2(n6337), .A3(n6338), .A4(n6339), .ZN(
        vectorData2[63]) );
  AOI22D1BWP U10829 ( .A1(n3569), .A2(\vrf/regTable[5][63] ), .B1(n3592), .B2(
        \vrf/regTable[7][63] ), .ZN(n6339) );
  AOI22D1BWP U10830 ( .A1(n3577), .A2(\vrf/regTable[4][63] ), .B1(n3591), .B2(
        \vrf/regTable[6][63] ), .ZN(n6338) );
  AOI22D1BWP U10831 ( .A1(n3571), .A2(\vrf/regTable[1][63] ), .B1(n3568), .B2(
        \vrf/regTable[3][63] ), .ZN(n6337) );
  AOI22D1BWP U10832 ( .A1(n3580), .A2(\vrf/regTable[0][63] ), .B1(n3566), .B2(
        \vrf/regTable[2][63] ), .ZN(n6336) );
  ND4D1BWP U10833 ( .A1(n6848), .A2(n6849), .A3(n6850), .A4(n6851), .ZN(
        vectorData2[191]) );
  AOI22D1BWP U10834 ( .A1(n3569), .A2(\vrf/regTable[5][191] ), .B1(n3578), 
        .B2(\vrf/regTable[7][191] ), .ZN(n6851) );
  AOI22D1BWP U10835 ( .A1(n3577), .A2(\vrf/regTable[4][191] ), .B1(n3573), 
        .B2(\vrf/regTable[6][191] ), .ZN(n6850) );
  AOI22D1BWP U10836 ( .A1(n3571), .A2(\vrf/regTable[1][191] ), .B1(n3597), 
        .B2(\vrf/regTable[3][191] ), .ZN(n6849) );
  AOI22D1BWP U10837 ( .A1(n3580), .A2(\vrf/regTable[0][191] ), .B1(n3593), 
        .B2(\vrf/regTable[2][191] ), .ZN(n6848) );
  AOI22D1BWP U10838 ( .A1(n5975), .A2(vectorData2[175]), .B1(n5984), .B2(
        vectorData2[223]), .ZN(n5889) );
  ND4D1BWP U10839 ( .A1(n6976), .A2(n6977), .A3(n6978), .A4(n6979), .ZN(
        vectorData2[223]) );
  AOI22D1BWP U10840 ( .A1(n3569), .A2(\vrf/regTable[5][223] ), .B1(n3592), 
        .B2(\vrf/regTable[7][223] ), .ZN(n6979) );
  AOI22D1BWP U10841 ( .A1(n3577), .A2(\vrf/regTable[4][223] ), .B1(n3591), 
        .B2(\vrf/regTable[6][223] ), .ZN(n6978) );
  AOI22D1BWP U10842 ( .A1(n3571), .A2(\vrf/regTable[1][223] ), .B1(n3568), 
        .B2(\vrf/regTable[3][223] ), .ZN(n6977) );
  AOI22D1BWP U10843 ( .A1(n3580), .A2(\vrf/regTable[0][223] ), .B1(n3566), 
        .B2(\vrf/regTable[2][223] ), .ZN(n6976) );
  ND4D1BWP U10844 ( .A1(n6784), .A2(n6785), .A3(n6786), .A4(n6787), .ZN(
        vectorData2[175]) );
  AOI22D1BWP U10845 ( .A1(n3569), .A2(\vrf/regTable[5][175] ), .B1(n3592), 
        .B2(\vrf/regTable[7][175] ), .ZN(n6787) );
  AOI22D1BWP U10846 ( .A1(n3577), .A2(\vrf/regTable[4][175] ), .B1(n3591), 
        .B2(\vrf/regTable[6][175] ), .ZN(n6786) );
  AOI22D1BWP U10847 ( .A1(n3571), .A2(\vrf/regTable[1][175] ), .B1(n3568), 
        .B2(\vrf/regTable[3][175] ), .ZN(n6785) );
  AOI22D1BWP U10848 ( .A1(n3580), .A2(\vrf/regTable[0][175] ), .B1(n3566), 
        .B2(\vrf/regTable[2][175] ), .ZN(n6784) );
  AOI22D1BWP U10849 ( .A1(n5977), .A2(vectorData2[143]), .B1(n5982), .B2(
        vectorData2[31]), .ZN(n5890) );
  ND4D1BWP U10850 ( .A1(n6208), .A2(n6209), .A3(n6210), .A4(n6211), .ZN(
        vectorData2[31]) );
  AOI22D1BWP U10851 ( .A1(n3569), .A2(\vrf/regTable[5][31] ), .B1(n3592), .B2(
        \vrf/regTable[7][31] ), .ZN(n6211) );
  AOI22D1BWP U10852 ( .A1(n3577), .A2(\vrf/regTable[4][31] ), .B1(n3591), .B2(
        \vrf/regTable[6][31] ), .ZN(n6210) );
  AOI22D1BWP U10853 ( .A1(n3571), .A2(\vrf/regTable[1][31] ), .B1(n3568), .B2(
        \vrf/regTable[3][31] ), .ZN(n6209) );
  AOI22D1BWP U10854 ( .A1(n3580), .A2(\vrf/regTable[0][31] ), .B1(n3566), .B2(
        \vrf/regTable[2][31] ), .ZN(n6208) );
  ND4D1BWP U10855 ( .A1(n6656), .A2(n6657), .A3(n6658), .A4(n6659), .ZN(
        vectorData2[143]) );
  AOI22D1BWP U10856 ( .A1(n3569), .A2(\vrf/regTable[5][143] ), .B1(n3592), 
        .B2(\vrf/regTable[7][143] ), .ZN(n6659) );
  AOI22D1BWP U10857 ( .A1(n3577), .A2(\vrf/regTable[4][143] ), .B1(n3591), 
        .B2(\vrf/regTable[6][143] ), .ZN(n6658) );
  AOI22D1BWP U10858 ( .A1(n3571), .A2(\vrf/regTable[1][143] ), .B1(n3568), 
        .B2(\vrf/regTable[3][143] ), .ZN(n6657) );
  AOI22D1BWP U10859 ( .A1(n3580), .A2(\vrf/regTable[0][143] ), .B1(n3566), 
        .B2(\vrf/regTable[2][143] ), .ZN(n6656) );
  AO222D1BWP U10860 ( .A1(scalarData2[8]), .A2(n4569), .B1(WR), .B2(n5971), 
        .C1(n4570), .C2(vectorData2[8]), .Z(dataOut[8]) );
  ND4D1BWP U10861 ( .A1(n6116), .A2(n6117), .A3(n6118), .A4(n6119), .ZN(
        vectorData2[8]) );
  AOI22D1BWP U10862 ( .A1(n3569), .A2(\vrf/regTable[5][8] ), .B1(n3578), .B2(
        \vrf/regTable[7][8] ), .ZN(n6119) );
  AOI22D1BWP U10863 ( .A1(n3577), .A2(\vrf/regTable[4][8] ), .B1(n3573), .B2(
        \vrf/regTable[6][8] ), .ZN(n6118) );
  AOI22D1BWP U10864 ( .A1(n3571), .A2(\vrf/regTable[1][8] ), .B1(n3597), .B2(
        \vrf/regTable[3][8] ), .ZN(n6117) );
  AOI22D1BWP U10865 ( .A1(n3580), .A2(\vrf/regTable[0][8] ), .B1(n3593), .B2(
        \vrf/regTable[2][8] ), .ZN(n6116) );
  ND3D1BWP U10866 ( .A1(n5970), .A2(n5969), .A3(n5968), .ZN(n5971) );
  AOI211XD0BWP U10867 ( .A1(n5977), .A2(vectorData2[136]), .B(n5967), .C(n5966), .ZN(n5968) );
  ND4D1BWP U10868 ( .A1(n5965), .A2(n5964), .A3(n5963), .A4(n5962), .ZN(n5966)
         );
  AOI22D1BWP U10869 ( .A1(n5981), .A2(vectorData2[184]), .B1(n5980), .B2(
        vectorData2[248]), .ZN(n5962) );
  ND4D1BWP U10870 ( .A1(n7076), .A2(n7077), .A3(n7078), .A4(n7079), .ZN(
        vectorData2[248]) );
  AOI22D1BWP U10871 ( .A1(n3569), .A2(\vrf/regTable[5][248] ), .B1(n3578), 
        .B2(\vrf/regTable[7][248] ), .ZN(n7079) );
  AOI22D1BWP U10872 ( .A1(n3577), .A2(\vrf/regTable[4][248] ), .B1(n3573), 
        .B2(\vrf/regTable[6][248] ), .ZN(n7078) );
  AOI22D1BWP U10873 ( .A1(n3571), .A2(\vrf/regTable[1][248] ), .B1(n3597), 
        .B2(\vrf/regTable[3][248] ), .ZN(n7077) );
  AOI22D1BWP U10874 ( .A1(n3580), .A2(\vrf/regTable[0][248] ), .B1(n3593), 
        .B2(\vrf/regTable[2][248] ), .ZN(n7076) );
  ND4D1BWP U10875 ( .A1(n6820), .A2(n6821), .A3(n6822), .A4(n6823), .ZN(
        vectorData2[184]) );
  AOI22D1BWP U10876 ( .A1(n3569), .A2(\vrf/regTable[5][184] ), .B1(n6083), 
        .B2(\vrf/regTable[7][184] ), .ZN(n6823) );
  AOI22D1BWP U10877 ( .A1(n3577), .A2(\vrf/regTable[4][184] ), .B1(n6081), 
        .B2(\vrf/regTable[6][184] ), .ZN(n6822) );
  AOI22D1BWP U10878 ( .A1(n3571), .A2(\vrf/regTable[1][184] ), .B1(n6079), 
        .B2(\vrf/regTable[3][184] ), .ZN(n6821) );
  AOI22D1BWP U10879 ( .A1(n3580), .A2(\vrf/regTable[0][184] ), .B1(n6075), 
        .B2(\vrf/regTable[2][184] ), .ZN(n6820) );
  AOI22D1BWP U10880 ( .A1(n5974), .A2(vectorData2[56]), .B1(n5972), .B2(
        vectorData2[120]), .ZN(n5963) );
  ND4D1BWP U10881 ( .A1(n6564), .A2(n6565), .A3(n6566), .A4(n6567), .ZN(
        vectorData2[120]) );
  AOI22D1BWP U10882 ( .A1(n3569), .A2(\vrf/regTable[5][120] ), .B1(n3578), 
        .B2(\vrf/regTable[7][120] ), .ZN(n6567) );
  AOI22D1BWP U10883 ( .A1(n3577), .A2(\vrf/regTable[4][120] ), .B1(n3573), 
        .B2(\vrf/regTable[6][120] ), .ZN(n6566) );
  AOI22D1BWP U10884 ( .A1(n3571), .A2(\vrf/regTable[1][120] ), .B1(n3597), 
        .B2(\vrf/regTable[3][120] ), .ZN(n6565) );
  AOI22D1BWP U10885 ( .A1(n3580), .A2(\vrf/regTable[0][120] ), .B1(n3593), 
        .B2(\vrf/regTable[2][120] ), .ZN(n6564) );
  ND4D1BWP U10886 ( .A1(n6308), .A2(n6309), .A3(n6310), .A4(n6311), .ZN(
        vectorData2[56]) );
  AOI22D1BWP U10887 ( .A1(n3569), .A2(\vrf/regTable[5][56] ), .B1(n3592), .B2(
        \vrf/regTable[7][56] ), .ZN(n6311) );
  AOI22D1BWP U10888 ( .A1(n3577), .A2(\vrf/regTable[4][56] ), .B1(n3591), .B2(
        \vrf/regTable[6][56] ), .ZN(n6310) );
  AOI22D1BWP U10889 ( .A1(n3571), .A2(\vrf/regTable[1][56] ), .B1(n3568), .B2(
        \vrf/regTable[3][56] ), .ZN(n6309) );
  AOI22D1BWP U10890 ( .A1(n3580), .A2(\vrf/regTable[0][56] ), .B1(n3566), .B2(
        \vrf/regTable[2][56] ), .ZN(n6308) );
  AOI22D1BWP U10891 ( .A1(n5979), .A2(vectorData2[88]), .B1(n5984), .B2(
        vectorData2[216]), .ZN(n5964) );
  ND4D1BWP U10892 ( .A1(n6948), .A2(n6949), .A3(n6950), .A4(n6951), .ZN(
        vectorData2[216]) );
  AOI22D1BWP U10893 ( .A1(n3569), .A2(\vrf/regTable[5][216] ), .B1(n3578), 
        .B2(\vrf/regTable[7][216] ), .ZN(n6951) );
  AOI22D1BWP U10894 ( .A1(n3577), .A2(\vrf/regTable[4][216] ), .B1(n3573), 
        .B2(\vrf/regTable[6][216] ), .ZN(n6950) );
  AOI22D1BWP U10895 ( .A1(n3571), .A2(\vrf/regTable[1][216] ), .B1(n3597), 
        .B2(\vrf/regTable[3][216] ), .ZN(n6949) );
  AOI22D1BWP U10896 ( .A1(n3580), .A2(\vrf/regTable[0][216] ), .B1(n3593), 
        .B2(\vrf/regTable[2][216] ), .ZN(n6948) );
  ND4D1BWP U10897 ( .A1(n6436), .A2(n6437), .A3(n6438), .A4(n6439), .ZN(
        vectorData2[88]) );
  AOI22D1BWP U10898 ( .A1(n6082), .A2(\vrf/regTable[5][88] ), .B1(n3592), .B2(
        \vrf/regTable[7][88] ), .ZN(n6439) );
  AOI22D1BWP U10899 ( .A1(n6080), .A2(\vrf/regTable[4][88] ), .B1(n3591), .B2(
        \vrf/regTable[6][88] ), .ZN(n6438) );
  AOI22D1BWP U10900 ( .A1(n6077), .A2(\vrf/regTable[1][88] ), .B1(n3568), .B2(
        \vrf/regTable[3][88] ), .ZN(n6437) );
  AOI22D1BWP U10901 ( .A1(n6073), .A2(\vrf/regTable[0][88] ), .B1(n3566), .B2(
        \vrf/regTable[2][88] ), .ZN(n6436) );
  AOI22D1BWP U10902 ( .A1(n5985), .A2(vectorData2[40]), .B1(n5982), .B2(
        vectorData2[24]), .ZN(n5965) );
  ND4D1BWP U10903 ( .A1(n6180), .A2(n6181), .A3(n6182), .A4(n6183), .ZN(
        vectorData2[24]) );
  AOI22D1BWP U10904 ( .A1(n3569), .A2(\vrf/regTable[5][24] ), .B1(n3592), .B2(
        \vrf/regTable[7][24] ), .ZN(n6183) );
  AOI22D1BWP U10905 ( .A1(n3577), .A2(\vrf/regTable[4][24] ), .B1(n3591), .B2(
        \vrf/regTable[6][24] ), .ZN(n6182) );
  AOI22D1BWP U10906 ( .A1(n3571), .A2(\vrf/regTable[1][24] ), .B1(n3568), .B2(
        \vrf/regTable[3][24] ), .ZN(n6181) );
  AOI22D1BWP U10907 ( .A1(n3580), .A2(\vrf/regTable[0][24] ), .B1(n3566), .B2(
        \vrf/regTable[2][24] ), .ZN(n6180) );
  ND4D1BWP U10908 ( .A1(n6244), .A2(n6245), .A3(n6246), .A4(n6247), .ZN(
        vectorData2[40]) );
  AOI22D1BWP U10909 ( .A1(n3569), .A2(\vrf/regTable[5][40] ), .B1(n3578), .B2(
        \vrf/regTable[7][40] ), .ZN(n6247) );
  AOI22D1BWP U10910 ( .A1(n3577), .A2(\vrf/regTable[4][40] ), .B1(n3573), .B2(
        \vrf/regTable[6][40] ), .ZN(n6246) );
  AOI22D1BWP U10911 ( .A1(n3571), .A2(\vrf/regTable[1][40] ), .B1(n3597), .B2(
        \vrf/regTable[3][40] ), .ZN(n6245) );
  AOI22D1BWP U10912 ( .A1(n3580), .A2(\vrf/regTable[0][40] ), .B1(n3593), .B2(
        \vrf/regTable[2][40] ), .ZN(n6244) );
  AO22D1BWP U10913 ( .A1(n5973), .A2(vectorData2[72]), .B1(n5983), .B2(
        vectorData2[152]), .Z(n5967) );
  ND4D1BWP U10914 ( .A1(n6692), .A2(n6693), .A3(n6694), .A4(n6695), .ZN(
        vectorData2[152]) );
  AOI22D1BWP U10915 ( .A1(n3569), .A2(\vrf/regTable[5][152] ), .B1(n3578), 
        .B2(\vrf/regTable[7][152] ), .ZN(n6695) );
  AOI22D1BWP U10916 ( .A1(n3577), .A2(\vrf/regTable[4][152] ), .B1(n3573), 
        .B2(\vrf/regTable[6][152] ), .ZN(n6694) );
  AOI22D1BWP U10917 ( .A1(n3571), .A2(\vrf/regTable[1][152] ), .B1(n3597), 
        .B2(\vrf/regTable[3][152] ), .ZN(n6693) );
  AOI22D1BWP U10918 ( .A1(n3580), .A2(\vrf/regTable[0][152] ), .B1(n3593), 
        .B2(\vrf/regTable[2][152] ), .ZN(n6692) );
  ND4D1BWP U10919 ( .A1(n6372), .A2(n6373), .A3(n6374), .A4(n6375), .ZN(
        vectorData2[72]) );
  AOI22D1BWP U10920 ( .A1(n3569), .A2(\vrf/regTable[5][72] ), .B1(n3578), .B2(
        \vrf/regTable[7][72] ), .ZN(n6375) );
  AOI22D1BWP U10921 ( .A1(n3577), .A2(\vrf/regTable[4][72] ), .B1(n3573), .B2(
        \vrf/regTable[6][72] ), .ZN(n6374) );
  AOI22D1BWP U10922 ( .A1(n3571), .A2(\vrf/regTable[1][72] ), .B1(n3597), .B2(
        \vrf/regTable[3][72] ), .ZN(n6373) );
  AOI22D1BWP U10923 ( .A1(n3580), .A2(\vrf/regTable[0][72] ), .B1(n3593), .B2(
        \vrf/regTable[2][72] ), .ZN(n6372) );
  ND4D1BWP U10924 ( .A1(n6628), .A2(n6629), .A3(n6630), .A4(n6631), .ZN(
        vectorData2[136]) );
  AOI22D1BWP U10925 ( .A1(n3569), .A2(\vrf/regTable[5][136] ), .B1(n3592), 
        .B2(\vrf/regTable[7][136] ), .ZN(n6631) );
  AOI22D1BWP U10926 ( .A1(n3577), .A2(\vrf/regTable[4][136] ), .B1(n3591), 
        .B2(\vrf/regTable[6][136] ), .ZN(n6630) );
  AOI22D1BWP U10927 ( .A1(n3571), .A2(\vrf/regTable[1][136] ), .B1(n3568), 
        .B2(\vrf/regTable[3][136] ), .ZN(n6629) );
  AOI22D1BWP U10928 ( .A1(n3580), .A2(\vrf/regTable[0][136] ), .B1(n3566), 
        .B2(\vrf/regTable[2][136] ), .ZN(n6628) );
  AOI22D1BWP U10929 ( .A1(n5975), .A2(vectorData2[168]), .B1(n5976), .B2(
        vectorData2[104]), .ZN(n5969) );
  ND4D1BWP U10930 ( .A1(n6500), .A2(n6501), .A3(n6502), .A4(n6503), .ZN(
        vectorData2[104]) );
  AOI22D1BWP U10931 ( .A1(n3569), .A2(\vrf/regTable[5][104] ), .B1(n3578), 
        .B2(\vrf/regTable[7][104] ), .ZN(n6503) );
  AOI22D1BWP U10932 ( .A1(n3577), .A2(\vrf/regTable[4][104] ), .B1(n3573), 
        .B2(\vrf/regTable[6][104] ), .ZN(n6502) );
  AOI22D1BWP U10933 ( .A1(n3571), .A2(\vrf/regTable[1][104] ), .B1(n3597), 
        .B2(\vrf/regTable[3][104] ), .ZN(n6501) );
  AOI22D1BWP U10934 ( .A1(n3580), .A2(\vrf/regTable[0][104] ), .B1(n3593), 
        .B2(\vrf/regTable[2][104] ), .ZN(n6500) );
  ND4D1BWP U10935 ( .A1(n6756), .A2(n6757), .A3(n6758), .A4(n6759), .ZN(
        vectorData2[168]) );
  AOI22D1BWP U10936 ( .A1(n3569), .A2(\vrf/regTable[5][168] ), .B1(n3578), 
        .B2(\vrf/regTable[7][168] ), .ZN(n6759) );
  AOI22D1BWP U10937 ( .A1(n3577), .A2(\vrf/regTable[4][168] ), .B1(n3573), 
        .B2(\vrf/regTable[6][168] ), .ZN(n6758) );
  AOI22D1BWP U10938 ( .A1(n3571), .A2(\vrf/regTable[1][168] ), .B1(n3597), 
        .B2(\vrf/regTable[3][168] ), .ZN(n6757) );
  AOI22D1BWP U10939 ( .A1(n3580), .A2(\vrf/regTable[0][168] ), .B1(n3593), 
        .B2(\vrf/regTable[2][168] ), .ZN(n6756) );
  AOI22D1BWP U10940 ( .A1(n5992), .A2(vectorData2[232]), .B1(n5978), .B2(
        vectorData2[200]), .ZN(n5970) );
  ND4D1BWP U10941 ( .A1(n6884), .A2(n6885), .A3(n6886), .A4(n6887), .ZN(
        vectorData2[200]) );
  AOI22D1BWP U10942 ( .A1(n3569), .A2(\vrf/regTable[5][200] ), .B1(n6083), 
        .B2(\vrf/regTable[7][200] ), .ZN(n6887) );
  AOI22D1BWP U10943 ( .A1(n3577), .A2(\vrf/regTable[4][200] ), .B1(n6081), 
        .B2(\vrf/regTable[6][200] ), .ZN(n6886) );
  AOI22D1BWP U10944 ( .A1(n3571), .A2(\vrf/regTable[1][200] ), .B1(n6079), 
        .B2(\vrf/regTable[3][200] ), .ZN(n6885) );
  AOI22D1BWP U10945 ( .A1(n3580), .A2(\vrf/regTable[0][200] ), .B1(n6075), 
        .B2(\vrf/regTable[2][200] ), .ZN(n6884) );
  ND4D1BWP U10946 ( .A1(n7012), .A2(n7013), .A3(n7014), .A4(n7015), .ZN(
        vectorData2[232]) );
  AOI22D1BWP U10947 ( .A1(n3569), .A2(\vrf/regTable[5][232] ), .B1(n3578), 
        .B2(\vrf/regTable[7][232] ), .ZN(n7015) );
  AOI22D1BWP U10948 ( .A1(n3577), .A2(\vrf/regTable[4][232] ), .B1(n3573), 
        .B2(\vrf/regTable[6][232] ), .ZN(n7014) );
  AOI22D1BWP U10949 ( .A1(n3571), .A2(\vrf/regTable[1][232] ), .B1(n3597), 
        .B2(\vrf/regTable[3][232] ), .ZN(n7013) );
  AOI22D1BWP U10950 ( .A1(n3580), .A2(\vrf/regTable[0][232] ), .B1(n3593), 
        .B2(\vrf/regTable[2][232] ), .ZN(n7012) );
  ND4D1BWP U10951 ( .A1(n8246), .A2(n8247), .A3(n8248), .A4(n8249), .ZN(
        scalarData2[8]) );
  AOI22D1BWP U10952 ( .A1(n8212), .A2(\srf/regTable[5][8] ), .B1(n8213), .B2(
        \srf/regTable[7][8] ), .ZN(n8249) );
  AOI22D1BWP U10953 ( .A1(n8210), .A2(\srf/regTable[4][8] ), .B1(n8211), .B2(
        \srf/regTable[6][8] ), .ZN(n8248) );
  AOI22D1BWP U10954 ( .A1(n8207), .A2(\srf/regTable[1][8] ), .B1(n8209), .B2(
        \srf/regTable[3][8] ), .ZN(n8247) );
  AOI22D1BWP U10955 ( .A1(n8203), .A2(\srf/regTable[0][8] ), .B1(n8205), .B2(
        \srf/regTable[2][8] ), .ZN(n8246) );
  AO222D1BWP U10956 ( .A1(WR), .A2(n5901), .B1(n4570), .B2(vectorData2[1]), 
        .C1(n4569), .C2(scalarData2[1]), .Z(dataOut[1]) );
  ND4D1BWP U10957 ( .A1(n8218), .A2(n8219), .A3(n8220), .A4(n8221), .ZN(
        scalarData2[1]) );
  AOI22D1BWP U10958 ( .A1(n8212), .A2(\srf/regTable[5][1] ), .B1(n8213), .B2(
        \srf/regTable[7][1] ), .ZN(n8221) );
  AOI22D1BWP U10959 ( .A1(n8210), .A2(\srf/regTable[4][1] ), .B1(n8211), .B2(
        \srf/regTable[6][1] ), .ZN(n8220) );
  AOI22D1BWP U10960 ( .A1(n8207), .A2(\srf/regTable[1][1] ), .B1(n8209), .B2(
        \srf/regTable[3][1] ), .ZN(n8219) );
  AOI22D1BWP U10961 ( .A1(n8203), .A2(\srf/regTable[0][1] ), .B1(n8205), .B2(
        \srf/regTable[2][1] ), .ZN(n8218) );
  ND4D1BWP U10962 ( .A1(n6088), .A2(n6089), .A3(n6090), .A4(n6091), .ZN(
        vectorData2[1]) );
  AOI22D1BWP U10963 ( .A1(n6082), .A2(\vrf/regTable[5][1] ), .B1(n3578), .B2(
        \vrf/regTable[7][1] ), .ZN(n6091) );
  AOI22D1BWP U10964 ( .A1(n3577), .A2(\vrf/regTable[4][1] ), .B1(n3573), .B2(
        \vrf/regTable[6][1] ), .ZN(n6090) );
  AOI22D1BWP U10965 ( .A1(n6077), .A2(\vrf/regTable[1][1] ), .B1(n3597), .B2(
        \vrf/regTable[3][1] ), .ZN(n6089) );
  AOI22D1BWP U10966 ( .A1(n3580), .A2(\vrf/regTable[0][1] ), .B1(n3593), .B2(
        \vrf/regTable[2][1] ), .ZN(n6088) );
  ND3D1BWP U10967 ( .A1(n5900), .A2(n5899), .A3(n5898), .ZN(n5901) );
  AOI211XD0BWP U10968 ( .A1(n5981), .A2(vectorData2[177]), .B(n5897), .C(n5896), .ZN(n5898) );
  ND4D1BWP U10969 ( .A1(n5895), .A2(n5894), .A3(n5893), .A4(n5892), .ZN(n5896)
         );
  AOI22D1BWP U10970 ( .A1(n5974), .A2(vectorData2[49]), .B1(n5980), .B2(
        vectorData2[241]), .ZN(n5892) );
  ND4D1BWP U10971 ( .A1(n7048), .A2(n7049), .A3(n7050), .A4(n7051), .ZN(
        vectorData2[241]) );
  AOI22D1BWP U10972 ( .A1(n3569), .A2(\vrf/regTable[5][241] ), .B1(n3592), 
        .B2(\vrf/regTable[7][241] ), .ZN(n7051) );
  AOI22D1BWP U10973 ( .A1(n3577), .A2(\vrf/regTable[4][241] ), .B1(n3591), 
        .B2(\vrf/regTable[6][241] ), .ZN(n7050) );
  AOI22D1BWP U10974 ( .A1(n3571), .A2(\vrf/regTable[1][241] ), .B1(n3568), 
        .B2(\vrf/regTable[3][241] ), .ZN(n7049) );
  AOI22D1BWP U10975 ( .A1(n3580), .A2(\vrf/regTable[0][241] ), .B1(n3566), 
        .B2(\vrf/regTable[2][241] ), .ZN(n7048) );
  ND4D1BWP U10976 ( .A1(n6280), .A2(n6281), .A3(n6282), .A4(n6283), .ZN(
        vectorData2[49]) );
  AOI22D1BWP U10977 ( .A1(n3569), .A2(\vrf/regTable[5][49] ), .B1(n3578), .B2(
        \vrf/regTable[7][49] ), .ZN(n6283) );
  AOI22D1BWP U10978 ( .A1(n3577), .A2(\vrf/regTable[4][49] ), .B1(n3573), .B2(
        \vrf/regTable[6][49] ), .ZN(n6282) );
  AOI22D1BWP U10979 ( .A1(n3571), .A2(\vrf/regTable[1][49] ), .B1(n3597), .B2(
        \vrf/regTable[3][49] ), .ZN(n6281) );
  AOI22D1BWP U10980 ( .A1(n3580), .A2(\vrf/regTable[0][49] ), .B1(n3593), .B2(
        \vrf/regTable[2][49] ), .ZN(n6280) );
  AOI22D1BWP U10981 ( .A1(n5979), .A2(vectorData2[81]), .B1(n5972), .B2(
        vectorData2[113]), .ZN(n5893) );
  ND4D1BWP U10982 ( .A1(n6536), .A2(n6537), .A3(n6538), .A4(n6539), .ZN(
        vectorData2[113]) );
  AOI22D1BWP U10983 ( .A1(n3569), .A2(\vrf/regTable[5][113] ), .B1(n3592), 
        .B2(\vrf/regTable[7][113] ), .ZN(n6539) );
  AOI22D1BWP U10984 ( .A1(n3577), .A2(\vrf/regTable[4][113] ), .B1(n3591), 
        .B2(\vrf/regTable[6][113] ), .ZN(n6538) );
  AOI22D1BWP U10985 ( .A1(n3571), .A2(\vrf/regTable[1][113] ), .B1(n3568), 
        .B2(\vrf/regTable[3][113] ), .ZN(n6537) );
  AOI22D1BWP U10986 ( .A1(n3580), .A2(\vrf/regTable[0][113] ), .B1(n3566), 
        .B2(\vrf/regTable[2][113] ), .ZN(n6536) );
  ND4D1BWP U10987 ( .A1(n6408), .A2(n6409), .A3(n6410), .A4(n6411), .ZN(
        vectorData2[81]) );
  AOI22D1BWP U10988 ( .A1(n3569), .A2(\vrf/regTable[5][81] ), .B1(n3592), .B2(
        \vrf/regTable[7][81] ), .ZN(n6411) );
  AOI22D1BWP U10989 ( .A1(n3577), .A2(\vrf/regTable[4][81] ), .B1(n3591), .B2(
        \vrf/regTable[6][81] ), .ZN(n6410) );
  AOI22D1BWP U10990 ( .A1(n3571), .A2(\vrf/regTable[1][81] ), .B1(n3568), .B2(
        \vrf/regTable[3][81] ), .ZN(n6409) );
  AOI22D1BWP U10991 ( .A1(n3580), .A2(\vrf/regTable[0][81] ), .B1(n3566), .B2(
        \vrf/regTable[2][81] ), .ZN(n6408) );
  AOI22D1BWP U10992 ( .A1(n5975), .A2(vectorData2[161]), .B1(n5984), .B2(
        vectorData2[209]), .ZN(n5894) );
  ND4D1BWP U10993 ( .A1(n6920), .A2(n6921), .A3(n6922), .A4(n6923), .ZN(
        vectorData2[209]) );
  AOI22D1BWP U10994 ( .A1(n3569), .A2(\vrf/regTable[5][209] ), .B1(n3592), 
        .B2(\vrf/regTable[7][209] ), .ZN(n6923) );
  AOI22D1BWP U10995 ( .A1(n3577), .A2(\vrf/regTable[4][209] ), .B1(n3591), 
        .B2(\vrf/regTable[6][209] ), .ZN(n6922) );
  AOI22D1BWP U10996 ( .A1(n3571), .A2(\vrf/regTable[1][209] ), .B1(n3568), 
        .B2(\vrf/regTable[3][209] ), .ZN(n6921) );
  AOI22D1BWP U10997 ( .A1(n3580), .A2(\vrf/regTable[0][209] ), .B1(n3566), 
        .B2(\vrf/regTable[2][209] ), .ZN(n6920) );
  ND4D1BWP U10998 ( .A1(n6728), .A2(n6729), .A3(n6730), .A4(n6731), .ZN(
        vectorData2[161]) );
  AOI22D1BWP U10999 ( .A1(n3569), .A2(\vrf/regTable[5][161] ), .B1(n3592), 
        .B2(\vrf/regTable[7][161] ), .ZN(n6731) );
  AOI22D1BWP U11000 ( .A1(n3577), .A2(\vrf/regTable[4][161] ), .B1(n3591), 
        .B2(\vrf/regTable[6][161] ), .ZN(n6730) );
  AOI22D1BWP U11001 ( .A1(n3571), .A2(\vrf/regTable[1][161] ), .B1(n3568), 
        .B2(\vrf/regTable[3][161] ), .ZN(n6729) );
  AOI22D1BWP U11002 ( .A1(n3580), .A2(\vrf/regTable[0][161] ), .B1(n3566), 
        .B2(\vrf/regTable[2][161] ), .ZN(n6728) );
  AOI22D1BWP U11003 ( .A1(n5978), .A2(vectorData2[193]), .B1(n5976), .B2(
        vectorData2[97]), .ZN(n5895) );
  ND4D1BWP U11004 ( .A1(n6472), .A2(n6473), .A3(n6474), .A4(n6475), .ZN(
        vectorData2[97]) );
  AOI22D1BWP U11005 ( .A1(n3569), .A2(\vrf/regTable[5][97] ), .B1(n3592), .B2(
        \vrf/regTable[7][97] ), .ZN(n6475) );
  AOI22D1BWP U11006 ( .A1(n3577), .A2(\vrf/regTable[4][97] ), .B1(n3591), .B2(
        \vrf/regTable[6][97] ), .ZN(n6474) );
  AOI22D1BWP U11007 ( .A1(n3571), .A2(\vrf/regTable[1][97] ), .B1(n3568), .B2(
        \vrf/regTable[3][97] ), .ZN(n6473) );
  AOI22D1BWP U11008 ( .A1(n3580), .A2(\vrf/regTable[0][97] ), .B1(n3566), .B2(
        \vrf/regTable[2][97] ), .ZN(n6472) );
  ND4D1BWP U11009 ( .A1(n6856), .A2(n6857), .A3(n6858), .A4(n6859), .ZN(
        vectorData2[193]) );
  AOI22D1BWP U11010 ( .A1(n3569), .A2(\vrf/regTable[5][193] ), .B1(n3578), 
        .B2(\vrf/regTable[7][193] ), .ZN(n6859) );
  AOI22D1BWP U11011 ( .A1(n3577), .A2(\vrf/regTable[4][193] ), .B1(n3573), 
        .B2(\vrf/regTable[6][193] ), .ZN(n6858) );
  AOI22D1BWP U11012 ( .A1(n3571), .A2(\vrf/regTable[1][193] ), .B1(n3597), 
        .B2(\vrf/regTable[3][193] ), .ZN(n6857) );
  AOI22D1BWP U11013 ( .A1(n3580), .A2(\vrf/regTable[0][193] ), .B1(n3593), 
        .B2(\vrf/regTable[2][193] ), .ZN(n6856) );
  AO22D1BWP U11014 ( .A1(n5985), .A2(vectorData2[33]), .B1(n5992), .B2(
        vectorData2[225]), .Z(n5897) );
  ND4D1BWP U11015 ( .A1(n6984), .A2(n6985), .A3(n6986), .A4(n6987), .ZN(
        vectorData2[225]) );
  AOI22D1BWP U11016 ( .A1(n3569), .A2(\vrf/regTable[5][225] ), .B1(n3578), 
        .B2(\vrf/regTable[7][225] ), .ZN(n6987) );
  AOI22D1BWP U11017 ( .A1(n3577), .A2(\vrf/regTable[4][225] ), .B1(n3573), 
        .B2(\vrf/regTable[6][225] ), .ZN(n6986) );
  AOI22D1BWP U11018 ( .A1(n3571), .A2(\vrf/regTable[1][225] ), .B1(n3597), 
        .B2(\vrf/regTable[3][225] ), .ZN(n6985) );
  AOI22D1BWP U11019 ( .A1(n3580), .A2(\vrf/regTable[0][225] ), .B1(n3593), 
        .B2(\vrf/regTable[2][225] ), .ZN(n6984) );
  ND4D1BWP U11020 ( .A1(n6216), .A2(n6217), .A3(n6218), .A4(n6219), .ZN(
        vectorData2[33]) );
  AOI22D1BWP U11021 ( .A1(n3569), .A2(\vrf/regTable[5][33] ), .B1(n3592), .B2(
        \vrf/regTable[7][33] ), .ZN(n6219) );
  AOI22D1BWP U11022 ( .A1(n3577), .A2(\vrf/regTable[4][33] ), .B1(n3591), .B2(
        \vrf/regTable[6][33] ), .ZN(n6218) );
  AOI22D1BWP U11023 ( .A1(n3571), .A2(\vrf/regTable[1][33] ), .B1(n3568), .B2(
        \vrf/regTable[3][33] ), .ZN(n6217) );
  AOI22D1BWP U11024 ( .A1(n3580), .A2(\vrf/regTable[0][33] ), .B1(n3566), .B2(
        \vrf/regTable[2][33] ), .ZN(n6216) );
  ND4D1BWP U11025 ( .A1(n6792), .A2(n6793), .A3(n6794), .A4(n6795), .ZN(
        vectorData2[177]) );
  AOI22D1BWP U11026 ( .A1(n3569), .A2(\vrf/regTable[5][177] ), .B1(n3592), 
        .B2(\vrf/regTable[7][177] ), .ZN(n6795) );
  AOI22D1BWP U11027 ( .A1(n3577), .A2(\vrf/regTable[4][177] ), .B1(n3591), 
        .B2(\vrf/regTable[6][177] ), .ZN(n6794) );
  AOI22D1BWP U11028 ( .A1(n3571), .A2(\vrf/regTable[1][177] ), .B1(n3568), 
        .B2(\vrf/regTable[3][177] ), .ZN(n6793) );
  AOI22D1BWP U11029 ( .A1(n3580), .A2(\vrf/regTable[0][177] ), .B1(n3566), 
        .B2(\vrf/regTable[2][177] ), .ZN(n6792) );
  AOI22D1BWP U11030 ( .A1(n5977), .A2(vectorData2[129]), .B1(n5973), .B2(
        vectorData2[65]), .ZN(n5899) );
  ND4D1BWP U11031 ( .A1(n6344), .A2(n6345), .A3(n6346), .A4(n6347), .ZN(
        vectorData2[65]) );
  AOI22D1BWP U11032 ( .A1(n3569), .A2(\vrf/regTable[5][65] ), .B1(n3592), .B2(
        \vrf/regTable[7][65] ), .ZN(n6347) );
  AOI22D1BWP U11033 ( .A1(n3577), .A2(\vrf/regTable[4][65] ), .B1(n3591), .B2(
        \vrf/regTable[6][65] ), .ZN(n6346) );
  AOI22D1BWP U11034 ( .A1(n3571), .A2(\vrf/regTable[1][65] ), .B1(n3568), .B2(
        \vrf/regTable[3][65] ), .ZN(n6345) );
  AOI22D1BWP U11035 ( .A1(n3580), .A2(\vrf/regTable[0][65] ), .B1(n3566), .B2(
        \vrf/regTable[2][65] ), .ZN(n6344) );
  ND4D1BWP U11036 ( .A1(n6600), .A2(n6601), .A3(n6602), .A4(n6603), .ZN(
        vectorData2[129]) );
  AOI22D1BWP U11037 ( .A1(n3569), .A2(\vrf/regTable[5][129] ), .B1(n3592), 
        .B2(\vrf/regTable[7][129] ), .ZN(n6603) );
  AOI22D1BWP U11038 ( .A1(n3577), .A2(\vrf/regTable[4][129] ), .B1(n3591), 
        .B2(\vrf/regTable[6][129] ), .ZN(n6602) );
  AOI22D1BWP U11039 ( .A1(n3571), .A2(\vrf/regTable[1][129] ), .B1(n3568), 
        .B2(\vrf/regTable[3][129] ), .ZN(n6601) );
  AOI22D1BWP U11040 ( .A1(n3580), .A2(\vrf/regTable[0][129] ), .B1(n3566), 
        .B2(\vrf/regTable[2][129] ), .ZN(n6600) );
  AOI22D1BWP U11041 ( .A1(n5983), .A2(vectorData2[145]), .B1(n5982), .B2(
        vectorData2[17]), .ZN(n5900) );
  ND4D1BWP U11042 ( .A1(n6152), .A2(n6153), .A3(n6154), .A4(n6155), .ZN(
        vectorData2[17]) );
  AOI22D1BWP U11043 ( .A1(n3569), .A2(\vrf/regTable[5][17] ), .B1(n3578), .B2(
        \vrf/regTable[7][17] ), .ZN(n6155) );
  AOI22D1BWP U11044 ( .A1(n3577), .A2(\vrf/regTable[4][17] ), .B1(n3573), .B2(
        \vrf/regTable[6][17] ), .ZN(n6154) );
  AOI22D1BWP U11045 ( .A1(n3571), .A2(\vrf/regTable[1][17] ), .B1(n3597), .B2(
        \vrf/regTable[3][17] ), .ZN(n6153) );
  AOI22D1BWP U11046 ( .A1(n3580), .A2(\vrf/regTable[0][17] ), .B1(n3593), .B2(
        \vrf/regTable[2][17] ), .ZN(n6152) );
  ND4D1BWP U11047 ( .A1(n6664), .A2(n6665), .A3(n6666), .A4(n6667), .ZN(
        vectorData2[145]) );
  AOI22D1BWP U11048 ( .A1(n3569), .A2(\vrf/regTable[5][145] ), .B1(n3578), 
        .B2(\vrf/regTable[7][145] ), .ZN(n6667) );
  AOI22D1BWP U11049 ( .A1(n3577), .A2(\vrf/regTable[4][145] ), .B1(n3573), 
        .B2(\vrf/regTable[6][145] ), .ZN(n6666) );
  AOI22D1BWP U11050 ( .A1(n3571), .A2(\vrf/regTable[1][145] ), .B1(n3597), 
        .B2(\vrf/regTable[3][145] ), .ZN(n6665) );
  AOI22D1BWP U11051 ( .A1(n3580), .A2(\vrf/regTable[0][145] ), .B1(n3593), 
        .B2(\vrf/regTable[2][145] ), .ZN(n6664) );
  AO222D1BWP U11052 ( .A1(scalarData2[10]), .A2(n4569), .B1(WR), .B2(n5841), 
        .C1(n4570), .C2(vectorData2[10]), .Z(dataOut[10]) );
  ND4D1BWP U11053 ( .A1(n6124), .A2(n6125), .A3(n6126), .A4(n6127), .ZN(
        vectorData2[10]) );
  AOI22D1BWP U11054 ( .A1(n3569), .A2(\vrf/regTable[5][10] ), .B1(n3592), .B2(
        \vrf/regTable[7][10] ), .ZN(n6127) );
  AOI22D1BWP U11055 ( .A1(n3577), .A2(\vrf/regTable[4][10] ), .B1(n3591), .B2(
        \vrf/regTable[6][10] ), .ZN(n6126) );
  AOI22D1BWP U11056 ( .A1(n3571), .A2(\vrf/regTable[1][10] ), .B1(n3568), .B2(
        \vrf/regTable[3][10] ), .ZN(n6125) );
  AOI22D1BWP U11057 ( .A1(n3580), .A2(\vrf/regTable[0][10] ), .B1(n3566), .B2(
        \vrf/regTable[2][10] ), .ZN(n6124) );
  ND3D1BWP U11058 ( .A1(n5840), .A2(n5839), .A3(n5838), .ZN(n5841) );
  AOI211XD0BWP U11059 ( .A1(n5985), .A2(vectorData2[42]), .B(n5837), .C(n5836), 
        .ZN(n5838) );
  ND4D1BWP U11060 ( .A1(n5835), .A2(n5834), .A3(n5833), .A4(n5832), .ZN(n5836)
         );
  AOI22D1BWP U11061 ( .A1(n5981), .A2(vectorData2[186]), .B1(n5977), .B2(
        vectorData2[138]), .ZN(n5832) );
  ND4D1BWP U11062 ( .A1(n6636), .A2(n6637), .A3(n6638), .A4(n6639), .ZN(
        vectorData2[138]) );
  AOI22D1BWP U11063 ( .A1(n3569), .A2(\vrf/regTable[5][138] ), .B1(n3592), 
        .B2(\vrf/regTable[7][138] ), .ZN(n6639) );
  AOI22D1BWP U11064 ( .A1(n3577), .A2(\vrf/regTable[4][138] ), .B1(n3591), 
        .B2(\vrf/regTable[6][138] ), .ZN(n6638) );
  AOI22D1BWP U11065 ( .A1(n3571), .A2(\vrf/regTable[1][138] ), .B1(n3568), 
        .B2(\vrf/regTable[3][138] ), .ZN(n6637) );
  AOI22D1BWP U11066 ( .A1(n3580), .A2(\vrf/regTable[0][138] ), .B1(n3566), 
        .B2(\vrf/regTable[2][138] ), .ZN(n6636) );
  ND4D1BWP U11067 ( .A1(n6828), .A2(n6829), .A3(n6830), .A4(n6831), .ZN(
        vectorData2[186]) );
  AOI22D1BWP U11068 ( .A1(n3569), .A2(\vrf/regTable[5][186] ), .B1(n3592), 
        .B2(\vrf/regTable[7][186] ), .ZN(n6831) );
  AOI22D1BWP U11069 ( .A1(n3577), .A2(\vrf/regTable[4][186] ), .B1(n3591), 
        .B2(\vrf/regTable[6][186] ), .ZN(n6830) );
  AOI22D1BWP U11070 ( .A1(n3571), .A2(\vrf/regTable[1][186] ), .B1(n3568), 
        .B2(\vrf/regTable[3][186] ), .ZN(n6829) );
  AOI22D1BWP U11071 ( .A1(n3580), .A2(\vrf/regTable[0][186] ), .B1(n3566), 
        .B2(\vrf/regTable[2][186] ), .ZN(n6828) );
  AOI22D1BWP U11072 ( .A1(n5992), .A2(vectorData2[234]), .B1(n5973), .B2(
        vectorData2[74]), .ZN(n5833) );
  ND4D1BWP U11073 ( .A1(n6380), .A2(n6381), .A3(n6382), .A4(n6383), .ZN(
        vectorData2[74]) );
  AOI22D1BWP U11074 ( .A1(n3569), .A2(\vrf/regTable[5][74] ), .B1(n3592), .B2(
        \vrf/regTable[7][74] ), .ZN(n6383) );
  AOI22D1BWP U11075 ( .A1(n3577), .A2(\vrf/regTable[4][74] ), .B1(n3591), .B2(
        \vrf/regTable[6][74] ), .ZN(n6382) );
  AOI22D1BWP U11076 ( .A1(n3571), .A2(\vrf/regTable[1][74] ), .B1(n3568), .B2(
        \vrf/regTable[3][74] ), .ZN(n6381) );
  AOI22D1BWP U11077 ( .A1(n3580), .A2(\vrf/regTable[0][74] ), .B1(n3566), .B2(
        \vrf/regTable[2][74] ), .ZN(n6380) );
  ND4D1BWP U11078 ( .A1(n7020), .A2(n7021), .A3(n7022), .A4(n7023), .ZN(
        vectorData2[234]) );
  AOI22D1BWP U11079 ( .A1(n3569), .A2(\vrf/regTable[5][234] ), .B1(n6083), 
        .B2(\vrf/regTable[7][234] ), .ZN(n7023) );
  AOI22D1BWP U11080 ( .A1(n3577), .A2(\vrf/regTable[4][234] ), .B1(n6081), 
        .B2(\vrf/regTable[6][234] ), .ZN(n7022) );
  AOI22D1BWP U11081 ( .A1(n3571), .A2(\vrf/regTable[1][234] ), .B1(n6079), 
        .B2(\vrf/regTable[3][234] ), .ZN(n7021) );
  AOI22D1BWP U11082 ( .A1(n3580), .A2(\vrf/regTable[0][234] ), .B1(n6075), 
        .B2(\vrf/regTable[2][234] ), .ZN(n7020) );
  AOI22D1BWP U11083 ( .A1(n5972), .A2(vectorData2[122]), .B1(n5980), .B2(
        vectorData2[250]), .ZN(n5834) );
  ND4D1BWP U11084 ( .A1(n7084), .A2(n7085), .A3(n7086), .A4(n7087), .ZN(
        vectorData2[250]) );
  AOI22D1BWP U11085 ( .A1(n3569), .A2(\vrf/regTable[5][250] ), .B1(n3578), 
        .B2(\vrf/regTable[7][250] ), .ZN(n7087) );
  AOI22D1BWP U11086 ( .A1(n3577), .A2(\vrf/regTable[4][250] ), .B1(n3573), 
        .B2(\vrf/regTable[6][250] ), .ZN(n7086) );
  AOI22D1BWP U11087 ( .A1(n3571), .A2(\vrf/regTable[1][250] ), .B1(n3597), 
        .B2(\vrf/regTable[3][250] ), .ZN(n7085) );
  AOI22D1BWP U11088 ( .A1(n3580), .A2(\vrf/regTable[0][250] ), .B1(n3593), 
        .B2(\vrf/regTable[2][250] ), .ZN(n7084) );
  ND4D1BWP U11089 ( .A1(n6572), .A2(n6573), .A3(n6574), .A4(n6575), .ZN(
        vectorData2[122]) );
  AOI22D1BWP U11090 ( .A1(n3569), .A2(\vrf/regTable[5][122] ), .B1(n3578), 
        .B2(\vrf/regTable[7][122] ), .ZN(n6575) );
  AOI22D1BWP U11091 ( .A1(n3577), .A2(\vrf/regTable[4][122] ), .B1(n3573), 
        .B2(\vrf/regTable[6][122] ), .ZN(n6574) );
  AOI22D1BWP U11092 ( .A1(n3571), .A2(\vrf/regTable[1][122] ), .B1(n3597), 
        .B2(\vrf/regTable[3][122] ), .ZN(n6573) );
  AOI22D1BWP U11093 ( .A1(n3580), .A2(\vrf/regTable[0][122] ), .B1(n3593), 
        .B2(\vrf/regTable[2][122] ), .ZN(n6572) );
  AOI22D1BWP U11094 ( .A1(n5974), .A2(vectorData2[58]), .B1(n5976), .B2(
        vectorData2[106]), .ZN(n5835) );
  ND4D1BWP U11095 ( .A1(n6508), .A2(n6509), .A3(n6510), .A4(n6511), .ZN(
        vectorData2[106]) );
  AOI22D1BWP U11096 ( .A1(n3569), .A2(\vrf/regTable[5][106] ), .B1(n3578), 
        .B2(\vrf/regTable[7][106] ), .ZN(n6511) );
  AOI22D1BWP U11097 ( .A1(n3577), .A2(\vrf/regTable[4][106] ), .B1(n3573), 
        .B2(\vrf/regTable[6][106] ), .ZN(n6510) );
  AOI22D1BWP U11098 ( .A1(n3571), .A2(\vrf/regTable[1][106] ), .B1(n3597), 
        .B2(\vrf/regTable[3][106] ), .ZN(n6509) );
  AOI22D1BWP U11099 ( .A1(n3580), .A2(\vrf/regTable[0][106] ), .B1(n3593), 
        .B2(\vrf/regTable[2][106] ), .ZN(n6508) );
  ND4D1BWP U11100 ( .A1(n6316), .A2(n6317), .A3(n6318), .A4(n6319), .ZN(
        vectorData2[58]) );
  AOI22D1BWP U11101 ( .A1(n3569), .A2(\vrf/regTable[5][58] ), .B1(n3592), .B2(
        \vrf/regTable[7][58] ), .ZN(n6319) );
  AOI22D1BWP U11102 ( .A1(n3577), .A2(\vrf/regTable[4][58] ), .B1(n3591), .B2(
        \vrf/regTable[6][58] ), .ZN(n6318) );
  AOI22D1BWP U11103 ( .A1(n3571), .A2(\vrf/regTable[1][58] ), .B1(n3568), .B2(
        \vrf/regTable[3][58] ), .ZN(n6317) );
  AOI22D1BWP U11104 ( .A1(n3580), .A2(\vrf/regTable[0][58] ), .B1(n3566), .B2(
        \vrf/regTable[2][58] ), .ZN(n6316) );
  AO22D1BWP U11105 ( .A1(n5979), .A2(vectorData2[90]), .B1(n5978), .B2(
        vectorData2[202]), .Z(n5837) );
  ND4D1BWP U11106 ( .A1(n6892), .A2(n6893), .A3(n6894), .A4(n6895), .ZN(
        vectorData2[202]) );
  AOI22D1BWP U11107 ( .A1(n3569), .A2(\vrf/regTable[5][202] ), .B1(n3578), 
        .B2(\vrf/regTable[7][202] ), .ZN(n6895) );
  AOI22D1BWP U11108 ( .A1(n3577), .A2(\vrf/regTable[4][202] ), .B1(n3573), 
        .B2(\vrf/regTable[6][202] ), .ZN(n6894) );
  AOI22D1BWP U11109 ( .A1(n3571), .A2(\vrf/regTable[1][202] ), .B1(n3597), 
        .B2(\vrf/regTable[3][202] ), .ZN(n6893) );
  AOI22D1BWP U11110 ( .A1(n3580), .A2(\vrf/regTable[0][202] ), .B1(n3593), 
        .B2(\vrf/regTable[2][202] ), .ZN(n6892) );
  ND4D1BWP U11111 ( .A1(n6444), .A2(n6445), .A3(n6446), .A4(n6447), .ZN(
        vectorData2[90]) );
  AOI22D1BWP U11112 ( .A1(n6082), .A2(\vrf/regTable[5][90] ), .B1(n3592), .B2(
        \vrf/regTable[7][90] ), .ZN(n6447) );
  AOI22D1BWP U11113 ( .A1(n6080), .A2(\vrf/regTable[4][90] ), .B1(n3591), .B2(
        \vrf/regTable[6][90] ), .ZN(n6446) );
  AOI22D1BWP U11114 ( .A1(n6077), .A2(\vrf/regTable[1][90] ), .B1(n3568), .B2(
        \vrf/regTable[3][90] ), .ZN(n6445) );
  AOI22D1BWP U11115 ( .A1(n6073), .A2(\vrf/regTable[0][90] ), .B1(n3566), .B2(
        \vrf/regTable[2][90] ), .ZN(n6444) );
  ND4D1BWP U11116 ( .A1(n6252), .A2(n6253), .A3(n6254), .A4(n6255), .ZN(
        vectorData2[42]) );
  AOI22D1BWP U11117 ( .A1(n3569), .A2(\vrf/regTable[5][42] ), .B1(n3578), .B2(
        \vrf/regTable[7][42] ), .ZN(n6255) );
  AOI22D1BWP U11118 ( .A1(n3577), .A2(\vrf/regTable[4][42] ), .B1(n3573), .B2(
        \vrf/regTable[6][42] ), .ZN(n6254) );
  AOI22D1BWP U11119 ( .A1(n3571), .A2(\vrf/regTable[1][42] ), .B1(n3597), .B2(
        \vrf/regTable[3][42] ), .ZN(n6253) );
  AOI22D1BWP U11120 ( .A1(n3580), .A2(\vrf/regTable[0][42] ), .B1(n3593), .B2(
        \vrf/regTable[2][42] ), .ZN(n6252) );
  AOI22D1BWP U11121 ( .A1(n5984), .A2(vectorData2[218]), .B1(n5983), .B2(
        vectorData2[154]), .ZN(n5839) );
  ND4D1BWP U11122 ( .A1(n6700), .A2(n6701), .A3(n6702), .A4(n6703), .ZN(
        vectorData2[154]) );
  AOI22D1BWP U11123 ( .A1(n3569), .A2(\vrf/regTable[5][154] ), .B1(n3592), 
        .B2(\vrf/regTable[7][154] ), .ZN(n6703) );
  AOI22D1BWP U11124 ( .A1(n3577), .A2(\vrf/regTable[4][154] ), .B1(n3591), 
        .B2(\vrf/regTable[6][154] ), .ZN(n6702) );
  AOI22D1BWP U11125 ( .A1(n3571), .A2(\vrf/regTable[1][154] ), .B1(n3568), 
        .B2(\vrf/regTable[3][154] ), .ZN(n6701) );
  AOI22D1BWP U11126 ( .A1(n3580), .A2(\vrf/regTable[0][154] ), .B1(n3566), 
        .B2(\vrf/regTable[2][154] ), .ZN(n6700) );
  ND4D1BWP U11127 ( .A1(n6956), .A2(n6957), .A3(n6958), .A4(n6959), .ZN(
        vectorData2[218]) );
  AOI22D1BWP U11128 ( .A1(n3569), .A2(\vrf/regTable[5][218] ), .B1(n3578), 
        .B2(\vrf/regTable[7][218] ), .ZN(n6959) );
  AOI22D1BWP U11129 ( .A1(n3577), .A2(\vrf/regTable[4][218] ), .B1(n3573), 
        .B2(\vrf/regTable[6][218] ), .ZN(n6958) );
  AOI22D1BWP U11130 ( .A1(n3571), .A2(\vrf/regTable[1][218] ), .B1(n3597), 
        .B2(\vrf/regTable[3][218] ), .ZN(n6957) );
  AOI22D1BWP U11131 ( .A1(n3580), .A2(\vrf/regTable[0][218] ), .B1(n3593), 
        .B2(\vrf/regTable[2][218] ), .ZN(n6956) );
  AOI22D1BWP U11132 ( .A1(n5975), .A2(vectorData2[170]), .B1(n5982), .B2(
        vectorData2[26]), .ZN(n5840) );
  ND4D1BWP U11133 ( .A1(n6188), .A2(n6189), .A3(n6190), .A4(n6191), .ZN(
        vectorData2[26]) );
  AOI22D1BWP U11134 ( .A1(n3569), .A2(\vrf/regTable[5][26] ), .B1(n3592), .B2(
        \vrf/regTable[7][26] ), .ZN(n6191) );
  AOI22D1BWP U11135 ( .A1(n6080), .A2(\vrf/regTable[4][26] ), .B1(n3591), .B2(
        \vrf/regTable[6][26] ), .ZN(n6190) );
  AOI22D1BWP U11136 ( .A1(n3571), .A2(\vrf/regTable[1][26] ), .B1(n3568), .B2(
        \vrf/regTable[3][26] ), .ZN(n6189) );
  AOI22D1BWP U11137 ( .A1(n6073), .A2(\vrf/regTable[0][26] ), .B1(n3566), .B2(
        \vrf/regTable[2][26] ), .ZN(n6188) );
  ND4D1BWP U11138 ( .A1(n6764), .A2(n6765), .A3(n6766), .A4(n6767), .ZN(
        vectorData2[170]) );
  AOI22D1BWP U11139 ( .A1(n3569), .A2(\vrf/regTable[5][170] ), .B1(n3578), 
        .B2(\vrf/regTable[7][170] ), .ZN(n6767) );
  AOI22D1BWP U11140 ( .A1(n3577), .A2(\vrf/regTable[4][170] ), .B1(n3573), 
        .B2(\vrf/regTable[6][170] ), .ZN(n6766) );
  AOI22D1BWP U11141 ( .A1(n3571), .A2(\vrf/regTable[1][170] ), .B1(n3597), 
        .B2(\vrf/regTable[3][170] ), .ZN(n6765) );
  AOI22D1BWP U11142 ( .A1(n3580), .A2(\vrf/regTable[0][170] ), .B1(n3593), 
        .B2(\vrf/regTable[2][170] ), .ZN(n6764) );
  ND4D1BWP U11143 ( .A1(n8254), .A2(n8255), .A3(n8256), .A4(n8257), .ZN(
        scalarData2[10]) );
  AOI22D1BWP U11144 ( .A1(n8212), .A2(\srf/regTable[5][10] ), .B1(n8213), .B2(
        \srf/regTable[7][10] ), .ZN(n8257) );
  AOI22D1BWP U11145 ( .A1(n8210), .A2(\srf/regTable[4][10] ), .B1(n8211), .B2(
        \srf/regTable[6][10] ), .ZN(n8256) );
  AOI22D1BWP U11146 ( .A1(n8207), .A2(\srf/regTable[1][10] ), .B1(n8209), .B2(
        \srf/regTable[3][10] ), .ZN(n8255) );
  AOI22D1BWP U11147 ( .A1(n8203), .A2(\srf/regTable[0][10] ), .B1(n8205), .B2(
        \srf/regTable[2][10] ), .ZN(n8254) );
  AO222D1BWP U11148 ( .A1(WR), .A2(n5851), .B1(n4570), .B2(vectorData2[11]), 
        .C1(n4569), .C2(scalarData2[11]), .Z(dataOut[11]) );
  ND4D1BWP U11149 ( .A1(n8258), .A2(n8259), .A3(n8260), .A4(n8261), .ZN(
        scalarData2[11]) );
  AOI22D1BWP U11150 ( .A1(n8212), .A2(\srf/regTable[5][11] ), .B1(n8213), .B2(
        \srf/regTable[7][11] ), .ZN(n8261) );
  AOI22D1BWP U11151 ( .A1(n8210), .A2(\srf/regTable[4][11] ), .B1(n8211), .B2(
        \srf/regTable[6][11] ), .ZN(n8260) );
  AOI22D1BWP U11152 ( .A1(n8207), .A2(\srf/regTable[1][11] ), .B1(n8209), .B2(
        \srf/regTable[3][11] ), .ZN(n8259) );
  AOI22D1BWP U11153 ( .A1(n8203), .A2(\srf/regTable[0][11] ), .B1(n8205), .B2(
        \srf/regTable[2][11] ), .ZN(n8258) );
  ND4D1BWP U11154 ( .A1(n6128), .A2(n6129), .A3(n6130), .A4(n6131), .ZN(
        vectorData2[11]) );
  AOI22D1BWP U11155 ( .A1(n3569), .A2(\vrf/regTable[5][11] ), .B1(n3592), .B2(
        \vrf/regTable[7][11] ), .ZN(n6131) );
  AOI22D1BWP U11156 ( .A1(n3577), .A2(\vrf/regTable[4][11] ), .B1(n3591), .B2(
        \vrf/regTable[6][11] ), .ZN(n6130) );
  AOI22D1BWP U11157 ( .A1(n3571), .A2(\vrf/regTable[1][11] ), .B1(n3568), .B2(
        \vrf/regTable[3][11] ), .ZN(n6129) );
  AOI22D1BWP U11158 ( .A1(n3580), .A2(\vrf/regTable[0][11] ), .B1(n3566), .B2(
        \vrf/regTable[2][11] ), .ZN(n6128) );
  ND3D1BWP U11159 ( .A1(n5850), .A2(n5849), .A3(n5848), .ZN(n5851) );
  AOI211XD0BWP U11160 ( .A1(n5978), .A2(vectorData2[203]), .B(n5847), .C(n5846), .ZN(n5848) );
  ND4D1BWP U11161 ( .A1(n5845), .A2(n5844), .A3(n5843), .A4(n5842), .ZN(n5846)
         );
  AOI22D1BWP U11162 ( .A1(n5979), .A2(vectorData2[91]), .B1(n5974), .B2(
        vectorData2[59]), .ZN(n5842) );
  ND4D1BWP U11163 ( .A1(n6320), .A2(n6321), .A3(n6322), .A4(n6323), .ZN(
        vectorData2[59]) );
  AOI22D1BWP U11164 ( .A1(n3569), .A2(\vrf/regTable[5][59] ), .B1(n3592), .B2(
        \vrf/regTable[7][59] ), .ZN(n6323) );
  AOI22D1BWP U11165 ( .A1(n3577), .A2(\vrf/regTable[4][59] ), .B1(n3591), .B2(
        \vrf/regTable[6][59] ), .ZN(n6322) );
  AOI22D1BWP U11166 ( .A1(n3571), .A2(\vrf/regTable[1][59] ), .B1(n3568), .B2(
        \vrf/regTable[3][59] ), .ZN(n6321) );
  AOI22D1BWP U11167 ( .A1(n3580), .A2(\vrf/regTable[0][59] ), .B1(n3566), .B2(
        \vrf/regTable[2][59] ), .ZN(n6320) );
  ND4D1BWP U11168 ( .A1(n6448), .A2(n6449), .A3(n6450), .A4(n6451), .ZN(
        vectorData2[91]) );
  AOI22D1BWP U11169 ( .A1(n3569), .A2(\vrf/regTable[5][91] ), .B1(n3592), .B2(
        \vrf/regTable[7][91] ), .ZN(n6451) );
  AOI22D1BWP U11170 ( .A1(n3577), .A2(\vrf/regTable[4][91] ), .B1(n3591), .B2(
        \vrf/regTable[6][91] ), .ZN(n6450) );
  AOI22D1BWP U11171 ( .A1(n3571), .A2(\vrf/regTable[1][91] ), .B1(n3568), .B2(
        \vrf/regTable[3][91] ), .ZN(n6449) );
  AOI22D1BWP U11172 ( .A1(n3580), .A2(\vrf/regTable[0][91] ), .B1(n3566), .B2(
        \vrf/regTable[2][91] ), .ZN(n6448) );
  AOI22D1BWP U11173 ( .A1(n5975), .A2(vectorData2[171]), .B1(n5982), .B2(
        vectorData2[27]), .ZN(n5843) );
  ND4D1BWP U11174 ( .A1(n6192), .A2(n6193), .A3(n6194), .A4(n6195), .ZN(
        vectorData2[27]) );
  AOI22D1BWP U11175 ( .A1(n3569), .A2(\vrf/regTable[5][27] ), .B1(n3578), .B2(
        \vrf/regTable[7][27] ), .ZN(n6195) );
  AOI22D1BWP U11176 ( .A1(n3577), .A2(\vrf/regTable[4][27] ), .B1(n3573), .B2(
        \vrf/regTable[6][27] ), .ZN(n6194) );
  AOI22D1BWP U11177 ( .A1(n3571), .A2(\vrf/regTable[1][27] ), .B1(n3597), .B2(
        \vrf/regTable[3][27] ), .ZN(n6193) );
  AOI22D1BWP U11178 ( .A1(n3580), .A2(\vrf/regTable[0][27] ), .B1(n3593), .B2(
        \vrf/regTable[2][27] ), .ZN(n6192) );
  ND4D1BWP U11179 ( .A1(n6768), .A2(n6769), .A3(n6770), .A4(n6771), .ZN(
        vectorData2[171]) );
  AOI22D1BWP U11180 ( .A1(n3569), .A2(\vrf/regTable[5][171] ), .B1(n3592), 
        .B2(\vrf/regTable[7][171] ), .ZN(n6771) );
  AOI22D1BWP U11181 ( .A1(n3577), .A2(\vrf/regTable[4][171] ), .B1(n3591), 
        .B2(\vrf/regTable[6][171] ), .ZN(n6770) );
  AOI22D1BWP U11182 ( .A1(n3571), .A2(\vrf/regTable[1][171] ), .B1(n3568), 
        .B2(\vrf/regTable[3][171] ), .ZN(n6769) );
  AOI22D1BWP U11183 ( .A1(n3580), .A2(\vrf/regTable[0][171] ), .B1(n3566), 
        .B2(\vrf/regTable[2][171] ), .ZN(n6768) );
  AOI22D1BWP U11184 ( .A1(n5981), .A2(vectorData2[187]), .B1(n5977), .B2(
        vectorData2[139]), .ZN(n5844) );
  ND4D1BWP U11185 ( .A1(n6640), .A2(n6641), .A3(n6642), .A4(n6643), .ZN(
        vectorData2[139]) );
  AOI22D1BWP U11186 ( .A1(n3569), .A2(\vrf/regTable[5][139] ), .B1(n3592), 
        .B2(\vrf/regTable[7][139] ), .ZN(n6643) );
  AOI22D1BWP U11187 ( .A1(n3577), .A2(\vrf/regTable[4][139] ), .B1(n3591), 
        .B2(\vrf/regTable[6][139] ), .ZN(n6642) );
  AOI22D1BWP U11188 ( .A1(n3571), .A2(\vrf/regTable[1][139] ), .B1(n3568), 
        .B2(\vrf/regTable[3][139] ), .ZN(n6641) );
  AOI22D1BWP U11189 ( .A1(n3580), .A2(\vrf/regTable[0][139] ), .B1(n3566), 
        .B2(\vrf/regTable[2][139] ), .ZN(n6640) );
  ND4D1BWP U11190 ( .A1(n6832), .A2(n6833), .A3(n6834), .A4(n6835), .ZN(
        vectorData2[187]) );
  AOI22D1BWP U11191 ( .A1(n3569), .A2(\vrf/regTable[5][187] ), .B1(n3592), 
        .B2(\vrf/regTable[7][187] ), .ZN(n6835) );
  AOI22D1BWP U11192 ( .A1(n3577), .A2(\vrf/regTable[4][187] ), .B1(n3591), 
        .B2(\vrf/regTable[6][187] ), .ZN(n6834) );
  AOI22D1BWP U11193 ( .A1(n3571), .A2(\vrf/regTable[1][187] ), .B1(n3568), 
        .B2(\vrf/regTable[3][187] ), .ZN(n6833) );
  AOI22D1BWP U11194 ( .A1(n3580), .A2(\vrf/regTable[0][187] ), .B1(n3566), 
        .B2(\vrf/regTable[2][187] ), .ZN(n6832) );
  AOI22D1BWP U11195 ( .A1(n5973), .A2(vectorData2[75]), .B1(n5976), .B2(
        vectorData2[107]), .ZN(n5845) );
  ND4D1BWP U11196 ( .A1(n6512), .A2(n6513), .A3(n6514), .A4(n6515), .ZN(
        vectorData2[107]) );
  AOI22D1BWP U11197 ( .A1(n3569), .A2(\vrf/regTable[5][107] ), .B1(n3578), 
        .B2(\vrf/regTable[7][107] ), .ZN(n6515) );
  AOI22D1BWP U11198 ( .A1(n3577), .A2(\vrf/regTable[4][107] ), .B1(n3573), 
        .B2(\vrf/regTable[6][107] ), .ZN(n6514) );
  AOI22D1BWP U11199 ( .A1(n3571), .A2(\vrf/regTable[1][107] ), .B1(n3597), 
        .B2(\vrf/regTable[3][107] ), .ZN(n6513) );
  AOI22D1BWP U11200 ( .A1(n3580), .A2(\vrf/regTable[0][107] ), .B1(n3593), 
        .B2(\vrf/regTable[2][107] ), .ZN(n6512) );
  ND4D1BWP U11201 ( .A1(n6384), .A2(n6385), .A3(n6386), .A4(n6387), .ZN(
        vectorData2[75]) );
  AOI22D1BWP U11202 ( .A1(n3569), .A2(\vrf/regTable[5][75] ), .B1(n3578), .B2(
        \vrf/regTable[7][75] ), .ZN(n6387) );
  AOI22D1BWP U11203 ( .A1(n3577), .A2(\vrf/regTable[4][75] ), .B1(n3573), .B2(
        \vrf/regTable[6][75] ), .ZN(n6386) );
  AOI22D1BWP U11204 ( .A1(n3571), .A2(\vrf/regTable[1][75] ), .B1(n3597), .B2(
        \vrf/regTable[3][75] ), .ZN(n6385) );
  AOI22D1BWP U11205 ( .A1(n3580), .A2(\vrf/regTable[0][75] ), .B1(n3593), .B2(
        \vrf/regTable[2][75] ), .ZN(n6384) );
  AO22D1BWP U11206 ( .A1(n5984), .A2(vectorData2[219]), .B1(n5980), .B2(
        vectorData2[251]), .Z(n5847) );
  ND4D1BWP U11207 ( .A1(n7088), .A2(n7089), .A3(n7090), .A4(n7091), .ZN(
        vectorData2[251]) );
  AOI22D1BWP U11208 ( .A1(n3569), .A2(\vrf/regTable[5][251] ), .B1(n6083), 
        .B2(\vrf/regTable[7][251] ), .ZN(n7091) );
  AOI22D1BWP U11209 ( .A1(n3577), .A2(\vrf/regTable[4][251] ), .B1(n6081), 
        .B2(\vrf/regTable[6][251] ), .ZN(n7090) );
  AOI22D1BWP U11210 ( .A1(n3571), .A2(\vrf/regTable[1][251] ), .B1(n6079), 
        .B2(\vrf/regTable[3][251] ), .ZN(n7089) );
  AOI22D1BWP U11211 ( .A1(n3580), .A2(\vrf/regTable[0][251] ), .B1(n6075), 
        .B2(\vrf/regTable[2][251] ), .ZN(n7088) );
  ND4D1BWP U11212 ( .A1(n6960), .A2(n6961), .A3(n6962), .A4(n6963), .ZN(
        vectorData2[219]) );
  AOI22D1BWP U11213 ( .A1(n3569), .A2(\vrf/regTable[5][219] ), .B1(n3592), 
        .B2(\vrf/regTable[7][219] ), .ZN(n6963) );
  AOI22D1BWP U11214 ( .A1(n3577), .A2(\vrf/regTable[4][219] ), .B1(n3591), 
        .B2(\vrf/regTable[6][219] ), .ZN(n6962) );
  AOI22D1BWP U11215 ( .A1(n3571), .A2(\vrf/regTable[1][219] ), .B1(n3568), 
        .B2(\vrf/regTable[3][219] ), .ZN(n6961) );
  AOI22D1BWP U11216 ( .A1(n3580), .A2(\vrf/regTable[0][219] ), .B1(n3566), 
        .B2(\vrf/regTable[2][219] ), .ZN(n6960) );
  ND4D1BWP U11217 ( .A1(n6896), .A2(n6897), .A3(n6898), .A4(n6899), .ZN(
        vectorData2[203]) );
  AOI22D1BWP U11218 ( .A1(n3569), .A2(\vrf/regTable[5][203] ), .B1(n3578), 
        .B2(\vrf/regTable[7][203] ), .ZN(n6899) );
  AOI22D1BWP U11219 ( .A1(n3577), .A2(\vrf/regTable[4][203] ), .B1(n3573), 
        .B2(\vrf/regTable[6][203] ), .ZN(n6898) );
  AOI22D1BWP U11220 ( .A1(n3571), .A2(\vrf/regTable[1][203] ), .B1(n3597), 
        .B2(\vrf/regTable[3][203] ), .ZN(n6897) );
  AOI22D1BWP U11221 ( .A1(n3580), .A2(\vrf/regTable[0][203] ), .B1(n3593), 
        .B2(\vrf/regTable[2][203] ), .ZN(n6896) );
  AOI22D1BWP U11222 ( .A1(n5985), .A2(vectorData2[43]), .B1(n5972), .B2(
        vectorData2[123]), .ZN(n5849) );
  ND4D1BWP U11223 ( .A1(n6576), .A2(n6577), .A3(n6578), .A4(n6579), .ZN(
        vectorData2[123]) );
  AOI22D1BWP U11224 ( .A1(n3569), .A2(\vrf/regTable[5][123] ), .B1(n3592), 
        .B2(\vrf/regTable[7][123] ), .ZN(n6579) );
  AOI22D1BWP U11225 ( .A1(n3577), .A2(\vrf/regTable[4][123] ), .B1(n3591), 
        .B2(\vrf/regTable[6][123] ), .ZN(n6578) );
  AOI22D1BWP U11226 ( .A1(n3571), .A2(\vrf/regTable[1][123] ), .B1(n3568), 
        .B2(\vrf/regTable[3][123] ), .ZN(n6577) );
  AOI22D1BWP U11227 ( .A1(n3580), .A2(\vrf/regTable[0][123] ), .B1(n3566), 
        .B2(\vrf/regTable[2][123] ), .ZN(n6576) );
  ND4D1BWP U11228 ( .A1(n6256), .A2(n6257), .A3(n6258), .A4(n6259), .ZN(
        vectorData2[43]) );
  AOI22D1BWP U11229 ( .A1(n3569), .A2(\vrf/regTable[5][43] ), .B1(n3578), .B2(
        \vrf/regTable[7][43] ), .ZN(n6259) );
  AOI22D1BWP U11230 ( .A1(n3577), .A2(\vrf/regTable[4][43] ), .B1(n3573), .B2(
        \vrf/regTable[6][43] ), .ZN(n6258) );
  AOI22D1BWP U11231 ( .A1(n3571), .A2(\vrf/regTable[1][43] ), .B1(n3597), .B2(
        \vrf/regTable[3][43] ), .ZN(n6257) );
  AOI22D1BWP U11232 ( .A1(n3580), .A2(\vrf/regTable[0][43] ), .B1(n3593), .B2(
        \vrf/regTable[2][43] ), .ZN(n6256) );
  AOI22D1BWP U11233 ( .A1(n5992), .A2(vectorData2[235]), .B1(n5983), .B2(
        vectorData2[155]), .ZN(n5850) );
  ND4D1BWP U11234 ( .A1(n6704), .A2(n6705), .A3(n6706), .A4(n6707), .ZN(
        vectorData2[155]) );
  AOI22D1BWP U11235 ( .A1(n3569), .A2(\vrf/regTable[5][155] ), .B1(n3578), 
        .B2(\vrf/regTable[7][155] ), .ZN(n6707) );
  AOI22D1BWP U11236 ( .A1(n3577), .A2(\vrf/regTable[4][155] ), .B1(n3573), 
        .B2(\vrf/regTable[6][155] ), .ZN(n6706) );
  AOI22D1BWP U11237 ( .A1(n3571), .A2(\vrf/regTable[1][155] ), .B1(n3597), 
        .B2(\vrf/regTable[3][155] ), .ZN(n6705) );
  AOI22D1BWP U11238 ( .A1(n3580), .A2(\vrf/regTable[0][155] ), .B1(n3593), 
        .B2(\vrf/regTable[2][155] ), .ZN(n6704) );
  ND4D1BWP U11239 ( .A1(n7024), .A2(n7025), .A3(n7026), .A4(n7027), .ZN(
        vectorData2[235]) );
  AOI22D1BWP U11240 ( .A1(n3569), .A2(\vrf/regTable[5][235] ), .B1(n3578), 
        .B2(\vrf/regTable[7][235] ), .ZN(n7027) );
  AOI22D1BWP U11241 ( .A1(n3577), .A2(\vrf/regTable[4][235] ), .B1(n3573), 
        .B2(\vrf/regTable[6][235] ), .ZN(n7026) );
  AOI22D1BWP U11242 ( .A1(n3571), .A2(\vrf/regTable[1][235] ), .B1(n3597), 
        .B2(\vrf/regTable[3][235] ), .ZN(n7025) );
  AOI22D1BWP U11243 ( .A1(n3580), .A2(\vrf/regTable[0][235] ), .B1(n3593), 
        .B2(\vrf/regTable[2][235] ), .ZN(n7024) );
  AO222D1BWP U11244 ( .A1(scalarData2[9]), .A2(n4569), .B1(WR), .B2(n5996), 
        .C1(n4570), .C2(vectorData2[9]), .Z(dataOut[9]) );
  ND4D1BWP U11245 ( .A1(n6120), .A2(n6121), .A3(n6122), .A4(n6123), .ZN(
        vectorData2[9]) );
  AOI22D1BWP U11246 ( .A1(n3569), .A2(\vrf/regTable[5][9] ), .B1(n3592), .B2(
        \vrf/regTable[7][9] ), .ZN(n6123) );
  AOI22D1BWP U11247 ( .A1(n3577), .A2(\vrf/regTable[4][9] ), .B1(n3591), .B2(
        \vrf/regTable[6][9] ), .ZN(n6122) );
  AOI22D1BWP U11248 ( .A1(n3571), .A2(\vrf/regTable[1][9] ), .B1(n3568), .B2(
        \vrf/regTable[3][9] ), .ZN(n6121) );
  AOI22D1BWP U11249 ( .A1(n3580), .A2(\vrf/regTable[0][9] ), .B1(n3566), .B2(
        \vrf/regTable[2][9] ), .ZN(n6120) );
  ND3D1BWP U11250 ( .A1(n5995), .A2(n5994), .A3(n5993), .ZN(n5996) );
  AOI211XD0BWP U11251 ( .A1(n5992), .A2(vectorData2[233]), .B(n5991), .C(n5990), .ZN(n5993) );
  ND4D1BWP U11252 ( .A1(n5989), .A2(n5988), .A3(n5987), .A4(n5986), .ZN(n5990)
         );
  AOI22D1BWP U11253 ( .A1(n5985), .A2(vectorData2[41]), .B1(n5984), .B2(
        vectorData2[217]), .ZN(n5986) );
  ND4D1BWP U11254 ( .A1(n6952), .A2(n6953), .A3(n6954), .A4(n6955), .ZN(
        vectorData2[217]) );
  AOI22D1BWP U11255 ( .A1(n3569), .A2(\vrf/regTable[5][217] ), .B1(n3578), 
        .B2(\vrf/regTable[7][217] ), .ZN(n6955) );
  AOI22D1BWP U11256 ( .A1(n3577), .A2(\vrf/regTable[4][217] ), .B1(n3573), 
        .B2(\vrf/regTable[6][217] ), .ZN(n6954) );
  AOI22D1BWP U11257 ( .A1(n3571), .A2(\vrf/regTable[1][217] ), .B1(n3597), 
        .B2(\vrf/regTable[3][217] ), .ZN(n6953) );
  AOI22D1BWP U11258 ( .A1(n3580), .A2(\vrf/regTable[0][217] ), .B1(n3593), 
        .B2(\vrf/regTable[2][217] ), .ZN(n6952) );
  ND4D1BWP U11259 ( .A1(n6248), .A2(n6249), .A3(n6250), .A4(n6251), .ZN(
        vectorData2[41]) );
  AOI22D1BWP U11260 ( .A1(n3569), .A2(\vrf/regTable[5][41] ), .B1(n3578), .B2(
        \vrf/regTable[7][41] ), .ZN(n6251) );
  AOI22D1BWP U11261 ( .A1(n3577), .A2(\vrf/regTable[4][41] ), .B1(n3573), .B2(
        \vrf/regTable[6][41] ), .ZN(n6250) );
  AOI22D1BWP U11262 ( .A1(n3571), .A2(\vrf/regTable[1][41] ), .B1(n3597), .B2(
        \vrf/regTable[3][41] ), .ZN(n6249) );
  AOI22D1BWP U11263 ( .A1(n3580), .A2(\vrf/regTable[0][41] ), .B1(n3593), .B2(
        \vrf/regTable[2][41] ), .ZN(n6248) );
  AOI22D1BWP U11264 ( .A1(n5983), .A2(vectorData2[153]), .B1(n5982), .B2(
        vectorData2[25]), .ZN(n5987) );
  ND4D1BWP U11265 ( .A1(n6184), .A2(n6185), .A3(n6186), .A4(n6187), .ZN(
        vectorData2[25]) );
  AOI22D1BWP U11266 ( .A1(n3569), .A2(\vrf/regTable[5][25] ), .B1(n3578), .B2(
        \vrf/regTable[7][25] ), .ZN(n6187) );
  AOI22D1BWP U11267 ( .A1(n3577), .A2(\vrf/regTable[4][25] ), .B1(n3573), .B2(
        \vrf/regTable[6][25] ), .ZN(n6186) );
  AOI22D1BWP U11268 ( .A1(n3571), .A2(\vrf/regTable[1][25] ), .B1(n3597), .B2(
        \vrf/regTable[3][25] ), .ZN(n6185) );
  AOI22D1BWP U11269 ( .A1(n3580), .A2(\vrf/regTable[0][25] ), .B1(n3593), .B2(
        \vrf/regTable[2][25] ), .ZN(n6184) );
  ND4D1BWP U11270 ( .A1(n6696), .A2(n6697), .A3(n6698), .A4(n6699), .ZN(
        vectorData2[153]) );
  AOI22D1BWP U11271 ( .A1(n3569), .A2(\vrf/regTable[5][153] ), .B1(n3578), 
        .B2(\vrf/regTable[7][153] ), .ZN(n6699) );
  AOI22D1BWP U11272 ( .A1(n3577), .A2(\vrf/regTable[4][153] ), .B1(n3573), 
        .B2(\vrf/regTable[6][153] ), .ZN(n6698) );
  AOI22D1BWP U11273 ( .A1(n3571), .A2(\vrf/regTable[1][153] ), .B1(n3597), 
        .B2(\vrf/regTable[3][153] ), .ZN(n6697) );
  AOI22D1BWP U11274 ( .A1(n3580), .A2(\vrf/regTable[0][153] ), .B1(n3593), 
        .B2(\vrf/regTable[2][153] ), .ZN(n6696) );
  AOI22D1BWP U11275 ( .A1(n5981), .A2(vectorData2[185]), .B1(n5980), .B2(
        vectorData2[249]), .ZN(n5988) );
  ND4D1BWP U11276 ( .A1(n7080), .A2(n7081), .A3(n7082), .A4(n7083), .ZN(
        vectorData2[249]) );
  AOI22D1BWP U11277 ( .A1(n3569), .A2(\vrf/regTable[5][249] ), .B1(n6083), 
        .B2(\vrf/regTable[7][249] ), .ZN(n7083) );
  AOI22D1BWP U11278 ( .A1(n3577), .A2(\vrf/regTable[4][249] ), .B1(n6081), 
        .B2(\vrf/regTable[6][249] ), .ZN(n7082) );
  AOI22D1BWP U11279 ( .A1(n3571), .A2(\vrf/regTable[1][249] ), .B1(n6079), 
        .B2(\vrf/regTable[3][249] ), .ZN(n7081) );
  AOI22D1BWP U11280 ( .A1(n3580), .A2(\vrf/regTable[0][249] ), .B1(n6075), 
        .B2(\vrf/regTable[2][249] ), .ZN(n7080) );
  ND4D1BWP U11281 ( .A1(n6824), .A2(n6825), .A3(n6826), .A4(n6827), .ZN(
        vectorData2[185]) );
  AOI22D1BWP U11282 ( .A1(n3569), .A2(\vrf/regTable[5][185] ), .B1(n3578), 
        .B2(\vrf/regTable[7][185] ), .ZN(n6827) );
  AOI22D1BWP U11283 ( .A1(n3577), .A2(\vrf/regTable[4][185] ), .B1(n3573), 
        .B2(\vrf/regTable[6][185] ), .ZN(n6826) );
  AOI22D1BWP U11284 ( .A1(n3571), .A2(\vrf/regTable[1][185] ), .B1(n3597), 
        .B2(\vrf/regTable[3][185] ), .ZN(n6825) );
  AOI22D1BWP U11285 ( .A1(n3580), .A2(\vrf/regTable[0][185] ), .B1(n3593), 
        .B2(\vrf/regTable[2][185] ), .ZN(n6824) );
  AOI22D1BWP U11286 ( .A1(n5979), .A2(vectorData2[89]), .B1(n5978), .B2(
        vectorData2[201]), .ZN(n5989) );
  ND4D1BWP U11287 ( .A1(n6888), .A2(n6889), .A3(n6890), .A4(n6891), .ZN(
        vectorData2[201]) );
  AOI22D1BWP U11288 ( .A1(n3569), .A2(\vrf/regTable[5][201] ), .B1(n3592), 
        .B2(\vrf/regTable[7][201] ), .ZN(n6891) );
  AOI22D1BWP U11289 ( .A1(n3577), .A2(\vrf/regTable[4][201] ), .B1(n3591), 
        .B2(\vrf/regTable[6][201] ), .ZN(n6890) );
  AOI22D1BWP U11290 ( .A1(n3571), .A2(\vrf/regTable[1][201] ), .B1(n3568), 
        .B2(\vrf/regTable[3][201] ), .ZN(n6889) );
  AOI22D1BWP U11291 ( .A1(n3580), .A2(\vrf/regTable[0][201] ), .B1(n3566), 
        .B2(\vrf/regTable[2][201] ), .ZN(n6888) );
  ND4D1BWP U11292 ( .A1(n6440), .A2(n6441), .A3(n6442), .A4(n6443), .ZN(
        vectorData2[89]) );
  AOI22D1BWP U11293 ( .A1(n6082), .A2(\vrf/regTable[5][89] ), .B1(n3592), .B2(
        \vrf/regTable[7][89] ), .ZN(n6443) );
  AOI22D1BWP U11294 ( .A1(n6080), .A2(\vrf/regTable[4][89] ), .B1(n3591), .B2(
        \vrf/regTable[6][89] ), .ZN(n6442) );
  AOI22D1BWP U11295 ( .A1(n6077), .A2(\vrf/regTable[1][89] ), .B1(n3568), .B2(
        \vrf/regTable[3][89] ), .ZN(n6441) );
  AOI22D1BWP U11296 ( .A1(n6073), .A2(\vrf/regTable[0][89] ), .B1(n3566), .B2(
        \vrf/regTable[2][89] ), .ZN(n6440) );
  AO22D1BWP U11297 ( .A1(n5977), .A2(vectorData2[137]), .B1(n5976), .B2(
        vectorData2[105]), .Z(n5991) );
  ND4D1BWP U11298 ( .A1(n6504), .A2(n6505), .A3(n6506), .A4(n6507), .ZN(
        vectorData2[105]) );
  AOI22D1BWP U11299 ( .A1(n3569), .A2(\vrf/regTable[5][105] ), .B1(n3578), 
        .B2(\vrf/regTable[7][105] ), .ZN(n6507) );
  AOI22D1BWP U11300 ( .A1(n3577), .A2(\vrf/regTable[4][105] ), .B1(n3573), 
        .B2(\vrf/regTable[6][105] ), .ZN(n6506) );
  AOI22D1BWP U11301 ( .A1(n3571), .A2(\vrf/regTable[1][105] ), .B1(n3597), 
        .B2(\vrf/regTable[3][105] ), .ZN(n6505) );
  AOI22D1BWP U11302 ( .A1(n3580), .A2(\vrf/regTable[0][105] ), .B1(n3593), 
        .B2(\vrf/regTable[2][105] ), .ZN(n6504) );
  ND4D1BWP U11303 ( .A1(n6632), .A2(n6633), .A3(n6634), .A4(n6635), .ZN(
        vectorData2[137]) );
  AOI22D1BWP U11304 ( .A1(n3569), .A2(\vrf/regTable[5][137] ), .B1(n3578), 
        .B2(\vrf/regTable[7][137] ), .ZN(n6635) );
  AOI22D1BWP U11305 ( .A1(n3577), .A2(\vrf/regTable[4][137] ), .B1(n3573), 
        .B2(\vrf/regTable[6][137] ), .ZN(n6634) );
  AOI22D1BWP U11306 ( .A1(n3571), .A2(\vrf/regTable[1][137] ), .B1(n3597), 
        .B2(\vrf/regTable[3][137] ), .ZN(n6633) );
  AOI22D1BWP U11307 ( .A1(n3580), .A2(\vrf/regTable[0][137] ), .B1(n3593), 
        .B2(\vrf/regTable[2][137] ), .ZN(n6632) );
  ND4D1BWP U11308 ( .A1(n7016), .A2(n7017), .A3(n7018), .A4(n7019), .ZN(
        vectorData2[233]) );
  AOI22D1BWP U11309 ( .A1(n3569), .A2(\vrf/regTable[5][233] ), .B1(n3578), 
        .B2(\vrf/regTable[7][233] ), .ZN(n7019) );
  AOI22D1BWP U11310 ( .A1(n3577), .A2(\vrf/regTable[4][233] ), .B1(n3573), 
        .B2(\vrf/regTable[6][233] ), .ZN(n7018) );
  AOI22D1BWP U11311 ( .A1(n3571), .A2(\vrf/regTable[1][233] ), .B1(n3597), 
        .B2(\vrf/regTable[3][233] ), .ZN(n7017) );
  AOI22D1BWP U11312 ( .A1(n3580), .A2(\vrf/regTable[0][233] ), .B1(n3593), 
        .B2(\vrf/regTable[2][233] ), .ZN(n7016) );
  AOI22D1BWP U11313 ( .A1(n5975), .A2(vectorData2[169]), .B1(n5974), .B2(
        vectorData2[57]), .ZN(n5994) );
  ND4D1BWP U11314 ( .A1(n6312), .A2(n6313), .A3(n6314), .A4(n6315), .ZN(
        vectorData2[57]) );
  AOI22D1BWP U11315 ( .A1(n3569), .A2(\vrf/regTable[5][57] ), .B1(n3592), .B2(
        \vrf/regTable[7][57] ), .ZN(n6315) );
  AOI22D1BWP U11316 ( .A1(n3577), .A2(\vrf/regTable[4][57] ), .B1(n3591), .B2(
        \vrf/regTable[6][57] ), .ZN(n6314) );
  AOI22D1BWP U11317 ( .A1(n3571), .A2(\vrf/regTable[1][57] ), .B1(n3568), .B2(
        \vrf/regTable[3][57] ), .ZN(n6313) );
  AOI22D1BWP U11318 ( .A1(n3580), .A2(\vrf/regTable[0][57] ), .B1(n3566), .B2(
        \vrf/regTable[2][57] ), .ZN(n6312) );
  ND4D1BWP U11319 ( .A1(n6760), .A2(n6761), .A3(n6762), .A4(n6763), .ZN(
        vectorData2[169]) );
  AOI22D1BWP U11320 ( .A1(n3569), .A2(\vrf/regTable[5][169] ), .B1(n3592), 
        .B2(\vrf/regTable[7][169] ), .ZN(n6763) );
  AOI22D1BWP U11321 ( .A1(n3577), .A2(\vrf/regTable[4][169] ), .B1(n3591), 
        .B2(\vrf/regTable[6][169] ), .ZN(n6762) );
  AOI22D1BWP U11322 ( .A1(n3571), .A2(\vrf/regTable[1][169] ), .B1(n3568), 
        .B2(\vrf/regTable[3][169] ), .ZN(n6761) );
  AOI22D1BWP U11323 ( .A1(n3580), .A2(\vrf/regTable[0][169] ), .B1(n3566), 
        .B2(\vrf/regTable[2][169] ), .ZN(n6760) );
  AOI22D1BWP U11324 ( .A1(n5973), .A2(vectorData2[73]), .B1(n5972), .B2(
        vectorData2[121]), .ZN(n5995) );
  ND4D1BWP U11325 ( .A1(n6568), .A2(n6569), .A3(n6570), .A4(n6571), .ZN(
        vectorData2[121]) );
  AOI22D1BWP U11326 ( .A1(n6082), .A2(\vrf/regTable[5][121] ), .B1(n3592), 
        .B2(\vrf/regTable[7][121] ), .ZN(n6571) );
  AOI22D1BWP U11327 ( .A1(n6080), .A2(\vrf/regTable[4][121] ), .B1(n3591), 
        .B2(\vrf/regTable[6][121] ), .ZN(n6570) );
  AOI22D1BWP U11328 ( .A1(n6077), .A2(\vrf/regTable[1][121] ), .B1(n3568), 
        .B2(\vrf/regTable[3][121] ), .ZN(n6569) );
  AOI22D1BWP U11329 ( .A1(n6073), .A2(\vrf/regTable[0][121] ), .B1(n3566), 
        .B2(\vrf/regTable[2][121] ), .ZN(n6568) );
  ND4D1BWP U11330 ( .A1(n6376), .A2(n6377), .A3(n6378), .A4(n6379), .ZN(
        vectorData2[73]) );
  AOI22D1BWP U11331 ( .A1(n3569), .A2(\vrf/regTable[5][73] ), .B1(n3578), .B2(
        \vrf/regTable[7][73] ), .ZN(n6379) );
  NR2XD0BWP U11332 ( .A1(n6076), .A2(n4622), .ZN(n6082) );
  AOI22D1BWP U11333 ( .A1(n3577), .A2(\vrf/regTable[4][73] ), .B1(n3573), .B2(
        \vrf/regTable[6][73] ), .ZN(n6378) );
  AOI22D1BWP U11334 ( .A1(n3571), .A2(\vrf/regTable[1][73] ), .B1(n3597), .B2(
        \vrf/regTable[3][73] ), .ZN(n6377) );
  NR2XD0BWP U11335 ( .A1(n6076), .A2(\vrf/N14 ), .ZN(n6077) );
  AOI22D1BWP U11336 ( .A1(n3580), .A2(\vrf/regTable[0][73] ), .B1(n3593), .B2(
        \vrf/regTable[2][73] ), .ZN(n6376) );
  NR2XD0BWP U11337 ( .A1(n5814), .A2(n5808), .ZN(n5985) );
  NR2XD0BWP U11338 ( .A1(n5810), .A2(n5816), .ZN(n5979) );
  NR2XD0BWP U11339 ( .A1(n5814), .A2(n5813), .ZN(n5976) );
  NR2XD0BWP U11340 ( .A1(n5810), .A2(n5814), .ZN(n5973) );
  NR2XD0BWP U11341 ( .A1(n5809), .A2(n5808), .ZN(n5975) );
  NR2XD0BWP U11342 ( .A1(n5809), .A2(n5813), .ZN(n5992) );
  NR2XD0BWP U11343 ( .A1(n5816), .A2(n5813), .ZN(n5972) );
  NR2XD0BWP U11344 ( .A1(n5810), .A2(n5815), .ZN(n5984) );
  NR2XD0BWP U11345 ( .A1(n5809), .A2(n5810), .ZN(n5978) );
  NR2XD0BWP U11346 ( .A1(n5809), .A2(n5805), .ZN(n5977) );
  NR2XD0BWP U11347 ( .A1(n5816), .A2(n5808), .ZN(n5974) );
  NR2XD0BWP U11348 ( .A1(n5815), .A2(n5808), .ZN(n5981) );
  NR2XD0BWP U11349 ( .A1(cycles[4]), .A2(n132), .ZN(n5806) );
  ND4D1BWP U11350 ( .A1(n8250), .A2(n8251), .A3(n8252), .A4(n8253), .ZN(
        scalarData2[9]) );
  AOI22D1BWP U11351 ( .A1(n8212), .A2(\srf/regTable[5][9] ), .B1(n8213), .B2(
        \srf/regTable[7][9] ), .ZN(n8253) );
  NR2XD0BWP U11352 ( .A1(n8208), .A2(n4622), .ZN(n8213) );
  NR2XD0BWP U11353 ( .A1(n8206), .A2(n4622), .ZN(n8212) );
  AOI22D1BWP U11354 ( .A1(n8210), .A2(\srf/regTable[4][9] ), .B1(n8211), .B2(
        \srf/regTable[6][9] ), .ZN(n8252) );
  NR2XD0BWP U11355 ( .A1(n8204), .A2(n4622), .ZN(n8211) );
  AOI22D1BWP U11356 ( .A1(n8207), .A2(\srf/regTable[1][9] ), .B1(n8209), .B2(
        \srf/regTable[3][9] ), .ZN(n8251) );
  NR2XD0BWP U11357 ( .A1(n8208), .A2(\vrf/N14 ), .ZN(n8209) );
  NR2XD0BWP U11358 ( .A1(n8206), .A2(\vrf/N14 ), .ZN(n8207) );
  AOI22D1BWP U11359 ( .A1(n8203), .A2(\srf/regTable[0][9] ), .B1(n8205), .B2(
        \srf/regTable[2][9] ), .ZN(n8250) );
  NR2XD0BWP U11360 ( .A1(n8204), .A2(\vrf/N14 ), .ZN(n8205) );
  OAI22D1BWP U11361 ( .A1(n153), .A2(n4551), .B1(n4553), .B2(n4555), .ZN(
        \vrf/N14 ) );
  IND3D1BWP U11362 ( .A1(Reset), .B1(n4392), .B2(n4616), .ZN(n3656) );
  IND2D1BWP U11363 ( .A1(Reset), .B1(n3717), .ZN(n3657) );
  ND3D1BWP U11364 ( .A1(n3714), .A2(n3715), .A3(n3713), .ZN(n4614) );
  AOI21D1BWP U11365 ( .A1(n4068), .A2(n3710), .B(n3709), .ZN(n3714) );
  AOI21D1BWP U11366 ( .A1(n3706), .A2(n3705), .B(Reset), .ZN(N152) );
  OAI21D1BWP U11367 ( .A1(code[0]), .A2(n3748), .B(n4553), .ZN(n3700) );
  ND3D1BWP U11368 ( .A1(n4394), .A2(n3716), .A3(n3563), .ZN(n3694) );
  OAI21D1BWP U11369 ( .A1(n3782), .A2(n3783), .B(n3682), .ZN(n3696) );
  ND3D1BWP U11370 ( .A1(n3562), .A2(n4394), .A3(n3719), .ZN(n3682) );
  OAI21D1BWP U11371 ( .A1(n3724), .A2(n3664), .B(n3723), .ZN(n3725) );
  ND3D1BWP U11372 ( .A1(n3663), .A2(n3563), .A3(n3612), .ZN(n3723) );
  ND3D1BWP U11373 ( .A1(n3562), .A2(state[1]), .A3(n3726), .ZN(n3724) );
  OAI21D1BWP U11374 ( .A1(n3787), .A2(n4554), .B(n3750), .ZN(n3718) );
  AN3XD1BWP U11375 ( .A1(n4394), .A2(n3681), .A3(n3563), .Z(n3660) );
  NR3D0BWP U11376 ( .A1(n3693), .A2(n3692), .A3(n3691), .ZN(n4573) );
  AOI31D1BWP U11377 ( .A1(n3690), .A2(n3689), .A3(n3699), .B(n4698), .ZN(n3691) );
  IND4D1BWP U11378 ( .A1(n3687), .B1(n3686), .B2(n3685), .B3(n4998), .ZN(n3693) );
  NR2XD0BWP U11379 ( .A1(n4552), .A2(n5812), .ZN(n3688) );
  AOI31D1BWP U11380 ( .A1(n3684), .A2(n3698), .A3(n3699), .B(n4392), .ZN(n4551) );
  OR2XD1BWP U11381 ( .A1(n4999), .A2(n5252), .Z(n3616) );
  INVD1BWP U11382 ( .I(n5334), .ZN(n4399) );
  AO22D1BWP U11383 ( .A1(n3652), .A2(n4718), .B1(n4717), .B2(n3678), .Z(n3618)
         );
  AO22D1BWP U11384 ( .A1(n3652), .A2(n4738), .B1(n4737), .B2(n3678), .Z(n3619)
         );
  NR2XD0BWP U11385 ( .A1(n4994), .A2(n4999), .ZN(n5187) );
  NR3D0BWP U11386 ( .A1(n3563), .A2(n4394), .A3(n4393), .ZN(n4060) );
  ND3D1BWP U11387 ( .A1(n6064), .A2(n6065), .A3(n6066), .ZN(result[10]) );
  FA1D0BWP U11388 ( .A(n4760), .B(n4759), .CI(n4758), .CO(n4757), .S(n4761) );
  FA1D0BWP U11389 ( .A(n4766), .B(n4765), .CI(n4764), .CO(n4763), .S(n4767) );
  FA1D0BWP U11390 ( .A(n4772), .B(n4771), .CI(n4770), .CO(n4769), .S(n4773) );
  FA1D0BWP U11391 ( .A(n4782), .B(n4781), .CI(n4780), .CO(n4779), .S(n4783) );
  NR3D0BWP U11392 ( .A1(\mult_x_153/n148 ), .A2(n4786), .A3(\mult_x_153/n136 ), 
        .ZN(\mult_x_153/n98 ) );
  MUX2ND0BWP U11393 ( .I0(n4612), .I1(n5793), .S(n4986), .ZN(\alu/N1019 ) );
  FA1D0BWP U11394 ( .A(op2[12]), .B(op1[12]), .CI(n4840), .CO(n4837), .S(
        \alu/N1016 ) );
  FA1D0BWP U11395 ( .A(op2[11]), .B(op1[11]), .CI(n4841), .CO(n4840), .S(
        \alu/N1015 ) );
  MUX2ND0BWP U11396 ( .I0(n5622), .I1(n3677), .S(n4842), .ZN(\alu/N1014 ) );
  MOAI22D0BWP U11397 ( .A1(n4874), .A2(n4866), .B1(n4635), .B2(n4875), .ZN(
        n4883) );
  NR3D0BWP U11398 ( .A1(n4881), .A2(n4922), .A3(n4965), .ZN(n4919) );
  FA1D0BWP U11399 ( .A(n4637), .B(n4884), .CI(n4883), .CO(n4885), .S(n4867) );
  MUX2ND0BWP U11400 ( .I0(result[4]), .I1(n4665), .S(n4971), .ZN(n4970) );
  MUX2ND0BWP U11401 ( .I0(result[15]), .I1(n6037), .S(n4984), .ZN(n4985) );
  NR4D0BWP U11402 ( .A1(result[5]), .A2(result[7]), .A3(result[8]), .A4(
        result[9]), .ZN(n4987) );
  INR3D0BWP U11403 ( .A1(n5208), .B1(n5207), .B2(n5240), .ZN(n5209) );
  INR3D0BWP U11404 ( .A1(n5221), .B1(n5220), .B2(n5240), .ZN(n5222) );
  INR3D0BWP U11405 ( .A1(n5242), .B1(n5241), .B2(n5240), .ZN(n5243) );
  FA1D0BWP U11406 ( .A(n5587), .B(n5586), .CI(n5585), .CO(n5588), .S(n5584) );
  FA1D0BWP U11407 ( .A(n5591), .B(n5590), .CI(n5589), .CO(n5598), .S(n5592) );
  FA1D0BWP U11408 ( .A(\mult_x_153/n30 ), .B(n5608), .CI(n5607), .CO(
        \intadd_33/B[9] ), .S(\intadd_33/B[8] ) );
  NR4D0BWP U11409 ( .A1(op1[1]), .A2(op1[9]), .A3(n5613), .A4(n5612), .ZN(
        n5621) );
  NR4D0BWP U11410 ( .A1(op1[2]), .A2(op1[0]), .A3(\alu/N87 ), .A4(n5614), .ZN(
        n5620) );
  NR4D0BWP U11411 ( .A1(op2[8]), .A2(op2[7]), .A3(op2[9]), .A4(op2[6]), .ZN(
        n5619) );
  NR4D0BWP U11412 ( .A1(op2[3]), .A2(op2[4]), .A3(\alu/N88 ), .A4(n5617), .ZN(
        n5618) );
  NR3D0BWP U11413 ( .A1(n4658), .A2(n5792), .A3(\alu/N683 ), .ZN(n5665) );
  MUX2ND0BWP U11414 ( .I0(n4658), .I1(\alu/N684 ), .S(n4657), .ZN(n5645) );
  MUX2ND0BWP U11415 ( .I0(\intadd_36/B[1] ), .I1(op1[12]), .S(n5642), .ZN(
        n5646) );
  MUX2ND0BWP U11416 ( .I0(n5655), .I1(n5647), .S(n5646), .ZN(n5657) );
  FA1D0BWP U11417 ( .A(n5650), .B(n5649), .CI(n5663), .CO(n5644), .S(n5669) );
  NR3D0BWP U11418 ( .A1(n5683), .A2(n5653), .A3(n5652), .ZN(n5691) );
  FA1D0BWP U11419 ( .A(n4660), .B(n5655), .CI(n5654), .CO(n5662), .S(n5661) );
  FA1D0BWP U11420 ( .A(n3653), .B(n5663), .CI(n5662), .CO(n5638), .S(n5664) );
  OA22D1BWP U11421 ( .A1(n4650), .A2(op2[15]), .B1(op1[15]), .B2(n5692), .Z(
        \alu/N634 ) );
  MOAI22D0BWP U11422 ( .A1(n5705), .A2(n4624), .B1(n4624), .B2(n5699), .ZN(
        n5700) );
  MUX2ND0BWP U11423 ( .I0(n5727), .I1(n5726), .S(n5739), .ZN(n5744) );
  MUX2ND0BWP U11424 ( .I0(n5736), .I1(n5728), .S(n5739), .ZN(n5741) );
  MUX2ND0BWP U11425 ( .I0(n5729), .I1(n5748), .S(n5739), .ZN(n5746) );
  MUX2ND0BWP U11426 ( .I0(n5785), .I1(n5784), .S(n5783), .ZN(n5791) );
  NR4D0BWP U11427 ( .A1(n5992), .A2(n5975), .A3(n5973), .A4(n5976), .ZN(n5830)
         );
  NR4D0BWP U11428 ( .A1(n5984), .A2(n5972), .A3(n5983), .A4(n5980), .ZN(n5829)
         );
  NR4D0BWP U11429 ( .A1(n5981), .A2(n5974), .A3(n5977), .A4(n5978), .ZN(n5828)
         );
endmodule
