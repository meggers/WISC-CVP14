module VectorRegFile ();

endmodule
