module DRAM_tb ();
  wire Clk1, Clk2;
  
  clock_source clocks(.Clk1(Clk1), .Clk2(Clk2));

endmodule
