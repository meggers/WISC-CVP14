module CVP14_tb();
  
endmodule
