module ScalarRegFile (rd_addr_1, rd_addr_2, wr_dst, wr_data, wr_en, data_1, data_2);

input rd_addr_1, rd_addr_2, wr_dst, wr_data, wr_en;
output data_1, data_2;



endmodule
