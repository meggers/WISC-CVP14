
module CVP14_DW01_addsub_0 ( A, B, CI, ADD_SUB, SUM, CO );
  input [4:0] A;
  input [4:0] B;
  output [4:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [5:0] carry;
  wire   [4:0] B_AS;
  assign carry[0] = ADD_SUB;

  XOR3D1BWP U1_4 ( .A1(A[4]), .A2(carry[0]), .A3(carry[4]), .Z(SUM[4]) );
  FA1D0BWP U1_3 ( .A(A[3]), .B(B_AS[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FA1D0BWP U1_2 ( .A(A[2]), .B(B_AS[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FA1D0BWP U1_1 ( .A(A[1]), .B(B_AS[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  FA1D0BWP U1_0 ( .A(A[0]), .B(B_AS[0]), .CI(carry[0]), .CO(carry[1]), .S(
        SUM[0]) );
  CKXOR2D0BWP U1 ( .A1(B[3]), .A2(carry[0]), .Z(B_AS[3]) );
  CKXOR2D0BWP U2 ( .A1(B[2]), .A2(carry[0]), .Z(B_AS[2]) );
  CKXOR2D0BWP U3 ( .A1(B[1]), .A2(carry[0]), .Z(B_AS[1]) );
  CKXOR2D0BWP U4 ( .A1(B[0]), .A2(carry[0]), .Z(B_AS[0]) );
endmodule


module CVP14_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [11:0] A;
  input [3:0] SH;
  output [11:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[3][11] , \ML_int[3][10] ,
         \ML_int[3][9] , \ML_int[3][8] , \ML_int[3][1] , \ML_int[3][0] ,
         \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] ,
         \ML_int[4][7] , \ML_int[4][6] , \ML_int[4][5] , \ML_int[4][4] ,
         \ML_int[4][3] , \ML_int[4][2] , n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14;
  assign B[11] = \ML_int[4][11] ;
  assign B[10] = \ML_int[4][10] ;
  assign B[9] = \ML_int[4][9] ;
  assign B[8] = \ML_int[4][8] ;
  assign B[7] = \ML_int[4][7] ;
  assign B[6] = \ML_int[4][6] ;
  assign B[5] = \ML_int[4][5] ;
  assign B[4] = \ML_int[4][4] ;
  assign B[3] = \ML_int[4][3] ;
  assign B[2] = \ML_int[4][2] ;

  MUX2D1BWP M1_3_11 ( .I0(\ML_int[3][11] ), .I1(n5), .S(SH[3]), .Z(
        \ML_int[4][11] ) );
  MUX2D1BWP M1_3_10 ( .I0(\ML_int[3][10] ), .I1(n6), .S(SH[3]), .Z(
        \ML_int[4][10] ) );
  MUX2D0BWP M1_2_9 ( .I0(\ML_int[2][9] ), .I1(\ML_int[2][5] ), .S(SH[2]), .Z(
        \ML_int[3][9] ) );
  MUX2D1BWP M1_3_9 ( .I0(\ML_int[3][9] ), .I1(\ML_int[3][1] ), .S(SH[3]), .Z(
        \ML_int[4][9] ) );
  MUX2D0BWP M1_2_8 ( .I0(\ML_int[2][8] ), .I1(\ML_int[2][4] ), .S(SH[2]), .Z(
        \ML_int[3][8] ) );
  MUX2D1BWP M1_3_8 ( .I0(\ML_int[3][8] ), .I1(\ML_int[3][0] ), .S(SH[3]), .Z(
        \ML_int[4][8] ) );
  MUX2D0BWP M1_0_1 ( .I0(A[1]), .I1(A[0]), .S(SH[0]), .Z(\ML_int[1][1] ) );
  MUX2D0BWP M1_0_9 ( .I0(A[9]), .I1(A[8]), .S(SH[0]), .Z(\ML_int[1][9] ) );
  MUX2D0BWP M1_0_5 ( .I0(A[5]), .I1(A[4]), .S(SH[0]), .Z(\ML_int[1][5] ) );
  MUX2D0BWP M1_0_6 ( .I0(A[6]), .I1(A[5]), .S(SH[0]), .Z(\ML_int[1][6] ) );
  MUX2D0BWP M1_0_2 ( .I0(A[2]), .I1(A[1]), .S(SH[0]), .Z(\ML_int[1][2] ) );
  MUX2D0BWP M1_0_11 ( .I0(A[11]), .I1(A[10]), .S(SH[0]), .Z(\ML_int[1][11] )
         );
  MUX2D0BWP M1_1_11 ( .I0(\ML_int[1][11] ), .I1(\ML_int[1][9] ), .S(SH[1]), 
        .Z(\ML_int[2][11] ) );
  MUX2D0BWP M1_2_11 ( .I0(\ML_int[2][11] ), .I1(\ML_int[2][7] ), .S(SH[2]), 
        .Z(\ML_int[3][11] ) );
  MUX2D0BWP M1_0_10 ( .I0(A[10]), .I1(A[9]), .S(SH[0]), .Z(\ML_int[1][10] ) );
  MUX2D0BWP M1_1_10 ( .I0(\ML_int[1][10] ), .I1(\ML_int[1][8] ), .S(SH[1]), 
        .Z(\ML_int[2][10] ) );
  MUX2D0BWP M1_2_10 ( .I0(\ML_int[2][10] ), .I1(\ML_int[2][6] ), .S(SH[2]), 
        .Z(\ML_int[3][10] ) );
  MUX2D0BWP M1_1_9 ( .I0(\ML_int[1][9] ), .I1(\ML_int[1][7] ), .S(SH[1]), .Z(
        \ML_int[2][9] ) );
  MUX2D0BWP M1_1_8 ( .I0(\ML_int[1][8] ), .I1(\ML_int[1][6] ), .S(SH[1]), .Z(
        \ML_int[2][8] ) );
  MUX2D0BWP M1_1_3 ( .I0(\ML_int[1][3] ), .I1(\ML_int[1][1] ), .S(SH[1]), .Z(
        \ML_int[2][3] ) );
  MUX2D0BWP M1_1_2 ( .I0(\ML_int[1][2] ), .I1(\ML_int[1][0] ), .S(SH[1]), .Z(
        \ML_int[2][2] ) );
  MUX2D0BWP M1_1_7 ( .I0(\ML_int[1][7] ), .I1(\ML_int[1][5] ), .S(SH[1]), .Z(
        \ML_int[2][7] ) );
  MUX2D0BWP M1_1_6 ( .I0(\ML_int[1][6] ), .I1(\ML_int[1][4] ), .S(SH[1]), .Z(
        \ML_int[2][6] ) );
  MUX2D0BWP M1_1_5 ( .I0(\ML_int[1][5] ), .I1(\ML_int[1][3] ), .S(SH[1]), .Z(
        \ML_int[2][5] ) );
  MUX2D0BWP M1_1_4 ( .I0(\ML_int[1][4] ), .I1(\ML_int[1][2] ), .S(SH[1]), .Z(
        \ML_int[2][4] ) );
  MUX2D0BWP M1_0_7 ( .I0(A[7]), .I1(A[6]), .S(SH[0]), .Z(\ML_int[1][7] ) );
  MUX2D0BWP M1_0_8 ( .I0(A[8]), .I1(A[7]), .S(SH[0]), .Z(\ML_int[1][8] ) );
  MUX2D0BWP M1_0_4 ( .I0(A[4]), .I1(A[3]), .S(SH[0]), .Z(\ML_int[1][4] ) );
  MUX2D0BWP M1_0_3 ( .I0(A[3]), .I1(A[2]), .S(SH[0]), .Z(\ML_int[1][3] ) );
  INR2D0BWP U3 ( .A1(A[0]), .B1(SH[0]), .ZN(\ML_int[1][0] ) );
  INVD1BWP U4 ( .I(SH[1]), .ZN(n10) );
  INVD1BWP U5 ( .I(n13), .ZN(n8) );
  INVD1BWP U6 ( .I(n14), .ZN(n9) );
  CKND0BWP U7 ( .I(SH[2]), .ZN(n7) );
  NR2XD0BWP U8 ( .A1(n1), .A2(SH[3]), .ZN(\ML_int[4][4] ) );
  MUX2ND0BWP U9 ( .I0(\ML_int[2][4] ), .I1(n9), .S(SH[2]), .ZN(n1) );
  NR2XD0BWP U10 ( .A1(n2), .A2(SH[3]), .ZN(\ML_int[4][5] ) );
  MUX2ND0BWP U11 ( .I0(\ML_int[2][5] ), .I1(n8), .S(SH[2]), .ZN(n2) );
  NR2XD0BWP U12 ( .A1(n3), .A2(SH[3]), .ZN(\ML_int[4][6] ) );
  MUX2ND0BWP U13 ( .I0(\ML_int[2][6] ), .I1(\ML_int[2][2] ), .S(SH[2]), .ZN(n3) );
  NR2XD0BWP U14 ( .A1(n4), .A2(SH[3]), .ZN(\ML_int[4][7] ) );
  MUX2ND0BWP U15 ( .I0(\ML_int[2][7] ), .I1(\ML_int[2][3] ), .S(SH[2]), .ZN(n4) );
  INVD1BWP U16 ( .I(n12), .ZN(n6) );
  INVD1BWP U17 ( .I(n11), .ZN(n5) );
  NR2D0BWP U18 ( .A1(n11), .A2(SH[3]), .ZN(\ML_int[4][3] ) );
  NR2D0BWP U19 ( .A1(n12), .A2(SH[3]), .ZN(\ML_int[4][2] ) );
  CKND2D0BWP U20 ( .A1(\ML_int[2][3] ), .A2(n7), .ZN(n11) );
  CKND2D0BWP U21 ( .A1(\ML_int[2][2] ), .A2(n7), .ZN(n12) );
  NR2D0BWP U22 ( .A1(SH[2]), .A2(n13), .ZN(\ML_int[3][1] ) );
  NR2D0BWP U23 ( .A1(SH[2]), .A2(n14), .ZN(\ML_int[3][0] ) );
  CKND2D0BWP U24 ( .A1(\ML_int[1][1] ), .A2(n10), .ZN(n13) );
  CKND2D0BWP U25 ( .A1(\ML_int[1][0] ), .A2(n10), .ZN(n14) );
endmodule


module CVP14_DW01_decode_0 ( A, B );
  input [4:0] A;
  output [31:0] B;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;

  INVD1BWP U2 ( .I(A[2]), .ZN(n3) );
  INVD1BWP U3 ( .I(A[0]), .ZN(n2) );
  INVD1BWP U4 ( .I(A[3]), .ZN(n1) );
  NR2D0BWP U5 ( .A1(n4), .A2(n5), .ZN(B[9]) );
  NR2D0BWP U6 ( .A1(n4), .A2(n6), .ZN(B[8]) );
  NR2D0BWP U7 ( .A1(n7), .A2(n8), .ZN(B[7]) );
  NR2D0BWP U8 ( .A1(n7), .A2(n9), .ZN(B[6]) );
  NR2D0BWP U9 ( .A1(n8), .A2(n10), .ZN(B[5]) );
  NR2D0BWP U10 ( .A1(n9), .A2(n10), .ZN(B[4]) );
  NR2D0BWP U11 ( .A1(n8), .A2(n11), .ZN(B[3]) );
  NR2D0BWP U12 ( .A1(n9), .A2(n11), .ZN(B[2]) );
  NR2D0BWP U13 ( .A1(n4), .A2(n8), .ZN(B[1]) );
  CKND2D0BWP U14 ( .A1(A[0]), .A2(n1), .ZN(n8) );
  NR2D0BWP U15 ( .A1(n6), .A2(n7), .ZN(B[14]) );
  CKND2D0BWP U16 ( .A1(A[1]), .A2(n12), .ZN(n7) );
  NR2D0BWP U17 ( .A1(n5), .A2(n10), .ZN(B[13]) );
  NR2D0BWP U18 ( .A1(n6), .A2(n10), .ZN(B[12]) );
  IND2D0BWP U19 ( .A1(A[1]), .B1(n12), .ZN(n10) );
  NR2D0BWP U20 ( .A1(n5), .A2(n11), .ZN(B[11]) );
  CKND2D0BWP U21 ( .A1(A[3]), .A2(A[0]), .ZN(n5) );
  NR2D0BWP U22 ( .A1(n6), .A2(n11), .ZN(B[10]) );
  IND3D0BWP U23 ( .A1(A[4]), .B1(n3), .B2(A[1]), .ZN(n11) );
  CKND2D0BWP U24 ( .A1(A[3]), .A2(n2), .ZN(n6) );
  NR2D0BWP U25 ( .A1(n4), .A2(n9), .ZN(B[0]) );
  CKND2D0BWP U26 ( .A1(n2), .A2(n1), .ZN(n9) );
  OR3D0BWP U27 ( .A1(n12), .A2(A[1]), .A3(A[4]), .Z(n4) );
  NR2D0BWP U28 ( .A1(n3), .A2(A[4]), .ZN(n12) );
endmodule


module CVP14_DW01_ash_1 ( A, DATA_TC, SH, SH_TC, B );
  input [255:0] A;
  input [8:0] SH;
  output [255:0] B;
  input DATA_TC, SH_TC;
  wire   \MR_int[4][1] , \MR_int[4][0] , \ML_int[4][14] , \ML_int[4][13] ,
         \ML_int[4][12] , \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] ,
         \ML_int[4][8] , \ML_int[4][7] , \ML_int[4][6] , \ML_int[4][5] ,
         \ML_int[4][4] , \ML_int[4][3] , \ML_int[4][2] , \ML_int[4][1] ,
         \ML_int[4][0] , \ML_int[5][32] , \ML_int[5][31] , \ML_int[5][30] ,
         \ML_int[5][29] , \ML_int[5][28] , \ML_int[5][27] , \ML_int[5][26] ,
         \ML_int[5][25] , \ML_int[5][24] , \ML_int[5][23] , \ML_int[5][22] ,
         \ML_int[5][21] , \ML_int[5][20] , \ML_int[5][19] , \ML_int[5][18] ,
         \ML_int[5][17] , \ML_int[5][16] , \ML_int[5][15] , \ML_int[5][14] ,
         \ML_int[5][13] , \ML_int[5][12] , \ML_int[5][11] , \ML_int[5][10] ,
         \ML_int[5][9] , \ML_int[5][8] , \ML_int[5][7] , \ML_int[5][6] ,
         \ML_int[5][5] , \ML_int[5][4] , \ML_int[5][3] , \ML_int[5][2] ,
         \ML_int[5][1] , \ML_int[5][0] , \ML_int[6][64] , \ML_int[6][63] ,
         \ML_int[6][62] , \ML_int[6][61] , \ML_int[6][60] , \ML_int[6][59] ,
         \ML_int[6][58] , \ML_int[6][57] , \ML_int[6][56] , \ML_int[6][55] ,
         \ML_int[6][54] , \ML_int[6][53] , \ML_int[6][52] , \ML_int[6][51] ,
         \ML_int[6][50] , \ML_int[6][49] , \ML_int[6][48] , \ML_int[6][47] ,
         \ML_int[6][46] , \ML_int[6][45] , \ML_int[6][44] , \ML_int[6][43] ,
         \ML_int[6][42] , \ML_int[6][41] , \ML_int[6][40] , \ML_int[6][39] ,
         \ML_int[6][38] , \ML_int[6][37] , \ML_int[6][36] , \ML_int[6][35] ,
         \ML_int[6][34] , \ML_int[6][33] , \ML_int[6][32] , \ML_int[6][31] ,
         \ML_int[6][30] , \ML_int[6][29] , \ML_int[6][28] , \ML_int[6][27] ,
         \ML_int[6][26] , \ML_int[6][25] , \ML_int[6][24] , \ML_int[6][23] ,
         \ML_int[6][22] , \ML_int[6][21] , \ML_int[6][20] , \ML_int[6][19] ,
         \ML_int[6][18] , \ML_int[6][17] , \ML_int[6][16] , \ML_int[6][15] ,
         \ML_int[6][14] , \ML_int[6][13] , \ML_int[6][12] , \ML_int[6][11] ,
         \ML_int[6][10] , \ML_int[6][9] , \ML_int[6][8] , \ML_int[6][7] ,
         \ML_int[6][6] , \ML_int[6][5] , \ML_int[6][4] , \ML_int[6][3] ,
         \ML_int[6][2] , \ML_int[6][1] , \ML_int[6][0] , \ML_int[7][128] ,
         \ML_int[7][127] , \ML_int[7][126] , \ML_int[7][125] ,
         \ML_int[7][124] , \ML_int[7][123] , \ML_int[7][122] ,
         \ML_int[7][121] , \ML_int[7][120] , \ML_int[7][119] ,
         \ML_int[7][118] , \ML_int[7][117] , \ML_int[7][116] ,
         \ML_int[7][115] , \ML_int[7][114] , \ML_int[7][113] ,
         \ML_int[7][112] , \ML_int[7][111] , \ML_int[7][110] ,
         \ML_int[7][109] , \ML_int[7][108] , \ML_int[7][107] ,
         \ML_int[7][106] , \ML_int[7][105] , \ML_int[7][104] ,
         \ML_int[7][103] , \ML_int[7][102] , \ML_int[7][101] ,
         \ML_int[7][100] , \ML_int[7][99] , \ML_int[7][98] , \ML_int[7][97] ,
         \ML_int[7][96] , \ML_int[7][95] , \ML_int[7][94] , \ML_int[7][93] ,
         \ML_int[7][92] , \ML_int[7][91] , \ML_int[7][90] , \ML_int[7][89] ,
         \ML_int[7][88] , \ML_int[7][87] , \ML_int[7][86] , \ML_int[7][85] ,
         \ML_int[7][84] , \ML_int[7][83] , \ML_int[7][82] , \ML_int[7][81] ,
         \ML_int[7][80] , \ML_int[7][79] , \ML_int[7][78] , \ML_int[7][77] ,
         \ML_int[7][76] , \ML_int[7][75] , \ML_int[7][74] , \ML_int[7][73] ,
         \ML_int[7][72] , \ML_int[7][71] , \ML_int[7][70] , \ML_int[7][69] ,
         \ML_int[7][68] , \ML_int[7][67] , \ML_int[7][66] , \ML_int[7][65] ,
         \ML_int[7][64] , \ML_int[8][255] , \ML_int[8][254] , \ML_int[8][253] ,
         \ML_int[8][252] , \ML_int[8][251] , \ML_int[8][250] ,
         \ML_int[8][249] , \ML_int[8][248] , \ML_int[8][247] ,
         \ML_int[8][246] , \ML_int[8][245] , \ML_int[8][244] ,
         \ML_int[8][243] , \ML_int[8][242] , \ML_int[8][241] ,
         \ML_int[8][240] , \ML_int[8][239] , \ML_int[8][238] ,
         \ML_int[8][237] , \ML_int[8][236] , \ML_int[8][235] ,
         \ML_int[8][234] , \ML_int[8][233] , \ML_int[8][232] ,
         \ML_int[8][231] , \ML_int[8][230] , \ML_int[8][229] ,
         \ML_int[8][228] , \ML_int[8][227] , \ML_int[8][226] ,
         \ML_int[8][225] , \ML_int[8][224] , \ML_int[8][223] ,
         \ML_int[8][222] , \ML_int[8][221] , \ML_int[8][220] ,
         \ML_int[8][219] , \ML_int[8][218] , \ML_int[8][217] ,
         \ML_int[8][216] , \ML_int[8][215] , \ML_int[8][214] ,
         \ML_int[8][213] , \ML_int[8][212] , \ML_int[8][211] ,
         \ML_int[8][210] , \ML_int[8][209] , \ML_int[8][208] ,
         \ML_int[8][207] , \ML_int[8][206] , \ML_int[8][205] ,
         \ML_int[8][204] , \ML_int[8][203] , \ML_int[8][202] ,
         \ML_int[8][201] , \ML_int[8][200] , \ML_int[8][199] ,
         \ML_int[8][198] , \ML_int[8][197] , \ML_int[8][196] ,
         \ML_int[8][195] , \ML_int[8][194] , \ML_int[8][193] ,
         \ML_int[8][192] , \ML_int[8][191] , \ML_int[8][190] ,
         \ML_int[8][189] , \ML_int[8][188] , \ML_int[8][187] ,
         \ML_int[8][186] , \ML_int[8][185] , \ML_int[8][184] ,
         \ML_int[8][183] , \ML_int[8][182] , \ML_int[8][181] ,
         \ML_int[8][180] , \ML_int[8][179] , \ML_int[8][178] ,
         \ML_int[8][177] , \ML_int[8][176] , \ML_int[8][175] ,
         \ML_int[8][174] , \ML_int[8][173] , \ML_int[8][172] ,
         \ML_int[8][171] , \ML_int[8][170] , \ML_int[8][169] ,
         \ML_int[8][168] , \ML_int[8][167] , \ML_int[8][166] ,
         \ML_int[8][165] , \ML_int[8][164] , \ML_int[8][163] ,
         \ML_int[8][162] , \ML_int[8][161] , \ML_int[8][160] ,
         \ML_int[8][159] , \ML_int[8][158] , \ML_int[8][157] ,
         \ML_int[8][156] , \ML_int[8][155] , \ML_int[8][154] ,
         \ML_int[8][153] , \ML_int[8][152] , \ML_int[8][151] ,
         \ML_int[8][150] , \ML_int[8][149] , \ML_int[8][148] ,
         \ML_int[8][147] , \ML_int[8][146] , \ML_int[8][145] ,
         \ML_int[8][144] , \ML_int[8][143] , \ML_int[8][142] ,
         \ML_int[8][141] , \ML_int[8][140] , \ML_int[8][139] ,
         \ML_int[8][138] , \ML_int[8][137] , \ML_int[8][136] ,
         \ML_int[8][135] , \ML_int[8][134] , \ML_int[8][133] ,
         \ML_int[8][132] , \ML_int[8][131] , \ML_int[8][130] ,
         \ML_int[8][129] , \ML_int[8][128] , \ML_int[9][255] ,
         \ML_int[9][254] , \ML_int[9][253] , \ML_int[9][252] ,
         \ML_int[9][251] , \ML_int[9][250] , \ML_int[9][249] ,
         \ML_int[9][248] , \ML_int[9][247] , \ML_int[9][246] ,
         \ML_int[9][245] , \ML_int[9][244] , \ML_int[9][243] ,
         \ML_int[9][242] , \ML_int[9][241] , \ML_int[9][240] ,
         \ML_int[9][239] , \ML_int[9][238] , \ML_int[9][237] ,
         \ML_int[9][236] , \ML_int[9][235] , \ML_int[9][234] ,
         \ML_int[9][233] , \ML_int[9][232] , \ML_int[9][231] ,
         \ML_int[9][230] , \ML_int[9][229] , \ML_int[9][228] ,
         \ML_int[9][227] , \ML_int[9][226] , \ML_int[9][225] ,
         \ML_int[9][224] , \ML_int[9][223] , \ML_int[9][222] ,
         \ML_int[9][221] , \ML_int[9][220] , \ML_int[9][219] ,
         \ML_int[9][218] , \ML_int[9][217] , \ML_int[9][216] ,
         \ML_int[9][215] , \ML_int[9][214] , \ML_int[9][213] ,
         \ML_int[9][212] , \ML_int[9][211] , \ML_int[9][210] ,
         \ML_int[9][209] , \ML_int[9][208] , \ML_int[9][207] ,
         \ML_int[9][206] , \ML_int[9][205] , \ML_int[9][204] ,
         \ML_int[9][203] , \ML_int[9][202] , \ML_int[9][201] ,
         \ML_int[9][200] , \ML_int[9][199] , \ML_int[9][198] ,
         \ML_int[9][197] , \ML_int[9][196] , \ML_int[9][195] ,
         \ML_int[9][194] , \ML_int[9][193] , \ML_int[9][192] ,
         \ML_int[9][191] , \ML_int[9][190] , \ML_int[9][189] ,
         \ML_int[9][188] , \ML_int[9][187] , \ML_int[9][186] ,
         \ML_int[9][185] , \ML_int[9][184] , \ML_int[9][183] ,
         \ML_int[9][182] , \ML_int[9][181] , \ML_int[9][180] ,
         \ML_int[9][179] , \ML_int[9][178] , \ML_int[9][177] ,
         \ML_int[9][176] , \ML_int[9][175] , \ML_int[9][174] ,
         \ML_int[9][173] , \ML_int[9][172] , \ML_int[9][171] ,
         \ML_int[9][170] , \ML_int[9][169] , \ML_int[9][168] ,
         \ML_int[9][167] , \ML_int[9][166] , \ML_int[9][165] ,
         \ML_int[9][164] , \ML_int[9][163] , \ML_int[9][162] ,
         \ML_int[9][161] , \ML_int[9][160] , \ML_int[9][159] ,
         \ML_int[9][158] , \ML_int[9][157] , \ML_int[9][156] ,
         \ML_int[9][155] , \ML_int[9][154] , \ML_int[9][153] ,
         \ML_int[9][152] , \ML_int[9][151] , \ML_int[9][150] ,
         \ML_int[9][149] , \ML_int[9][148] , \ML_int[9][147] ,
         \ML_int[9][146] , \ML_int[9][145] , \ML_int[9][144] ,
         \ML_int[9][143] , \ML_int[9][142] , \ML_int[9][141] ,
         \ML_int[9][140] , \ML_int[9][139] , \ML_int[9][138] ,
         \ML_int[9][137] , \ML_int[9][136] , \ML_int[9][135] ,
         \ML_int[9][134] , \ML_int[9][133] , \ML_int[9][132] ,
         \ML_int[9][131] , \ML_int[9][130] , \ML_int[9][129] ,
         \ML_int[9][128] , \ML_int[9][127] , \ML_int[9][126] ,
         \ML_int[9][125] , \ML_int[9][124] , \ML_int[9][123] ,
         \ML_int[9][122] , \ML_int[9][121] , \ML_int[9][120] ,
         \ML_int[9][119] , \ML_int[9][118] , \ML_int[9][117] ,
         \ML_int[9][116] , \ML_int[9][115] , \ML_int[9][114] ,
         \ML_int[9][113] , \ML_int[9][112] , \ML_int[9][111] ,
         \ML_int[9][110] , \ML_int[9][109] , \ML_int[9][108] ,
         \ML_int[9][107] , \ML_int[9][106] , \ML_int[9][105] ,
         \ML_int[9][104] , \ML_int[9][103] , \ML_int[9][102] ,
         \ML_int[9][101] , \ML_int[9][100] , \ML_int[9][99] , \ML_int[9][98] ,
         \ML_int[9][97] , \ML_int[9][96] , \ML_int[9][95] , \ML_int[9][94] ,
         \ML_int[9][93] , \ML_int[9][92] , \ML_int[9][91] , \ML_int[9][90] ,
         \ML_int[9][89] , \ML_int[9][88] , \ML_int[9][87] , \ML_int[9][86] ,
         \ML_int[9][85] , \ML_int[9][84] , \ML_int[9][83] , \ML_int[9][82] ,
         \ML_int[9][81] , \ML_int[9][80] , \ML_int[9][79] , \ML_int[9][78] ,
         \ML_int[9][77] , \ML_int[9][76] , \ML_int[9][75] , \ML_int[9][74] ,
         \ML_int[9][73] , \ML_int[9][72] , \ML_int[9][71] , \ML_int[9][70] ,
         \ML_int[9][69] , \ML_int[9][68] , \ML_int[9][67] , \ML_int[9][66] ,
         \ML_int[9][65] , \ML_int[9][64] , \ML_int[9][63] , \ML_int[9][62] ,
         \ML_int[9][61] , \ML_int[9][60] , \ML_int[9][59] , \ML_int[9][58] ,
         \ML_int[9][57] , \ML_int[9][56] , \ML_int[9][55] , \ML_int[9][54] ,
         \ML_int[9][53] , \ML_int[9][52] , \ML_int[9][51] , \ML_int[9][50] ,
         \ML_int[9][49] , \ML_int[9][48] , \ML_int[9][47] , \ML_int[9][46] ,
         \ML_int[9][45] , \ML_int[9][44] , \ML_int[9][43] , \ML_int[9][42] ,
         \ML_int[9][41] , \ML_int[9][40] , \ML_int[9][39] , \ML_int[9][38] ,
         \ML_int[9][37] , \ML_int[9][36] , \ML_int[9][35] , \ML_int[9][34] ,
         \ML_int[9][33] , \ML_int[9][32] , \ML_int[9][31] , \ML_int[9][30] ,
         \ML_int[9][29] , \ML_int[9][28] , \ML_int[9][27] , \ML_int[9][26] ,
         \ML_int[9][25] , \ML_int[9][24] , \ML_int[9][23] , \ML_int[9][22] ,
         \ML_int[9][21] , \ML_int[9][20] , \ML_int[9][19] , \ML_int[9][18] ,
         \ML_int[9][17] , \ML_int[9][16] , \ML_int[9][15] , \ML_int[9][14] ,
         \ML_int[9][13] , \ML_int[9][12] , \ML_int[9][11] , \ML_int[9][10] ,
         \ML_int[9][9] , \ML_int[9][8] , \ML_int[9][7] , \ML_int[9][6] ,
         \ML_int[9][5] , \ML_int[9][4] , \ML_int[9][3] , \ML_int[9][2] ,
         \ML_int[9][1] , \ML_int[9][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155;
  assign \MR_int[4][1]  = A[16];
  assign \MR_int[4][0]  = A[15];
  assign \ML_int[4][14]  = A[14];
  assign \ML_int[4][13]  = A[13];
  assign \ML_int[4][12]  = A[12];
  assign \ML_int[4][11]  = A[11];
  assign \ML_int[4][10]  = A[10];
  assign \ML_int[4][9]  = A[9];
  assign \ML_int[4][8]  = A[8];
  assign \ML_int[4][7]  = A[7];
  assign \ML_int[4][6]  = A[6];
  assign \ML_int[4][5]  = A[5];
  assign \ML_int[4][4]  = A[4];
  assign \ML_int[4][3]  = A[3];
  assign \ML_int[4][2]  = A[2];
  assign \ML_int[4][1]  = A[1];
  assign \ML_int[4][0]  = A[0];
  assign B[255] = \ML_int[9][255] ;
  assign B[254] = \ML_int[9][254] ;
  assign B[253] = \ML_int[9][253] ;
  assign B[252] = \ML_int[9][252] ;
  assign B[251] = \ML_int[9][251] ;
  assign B[250] = \ML_int[9][250] ;
  assign B[249] = \ML_int[9][249] ;
  assign B[248] = \ML_int[9][248] ;
  assign B[247] = \ML_int[9][247] ;
  assign B[246] = \ML_int[9][246] ;
  assign B[245] = \ML_int[9][245] ;
  assign B[244] = \ML_int[9][244] ;
  assign B[243] = \ML_int[9][243] ;
  assign B[242] = \ML_int[9][242] ;
  assign B[241] = \ML_int[9][241] ;
  assign B[240] = \ML_int[9][240] ;
  assign B[239] = \ML_int[9][239] ;
  assign B[238] = \ML_int[9][238] ;
  assign B[237] = \ML_int[9][237] ;
  assign B[236] = \ML_int[9][236] ;
  assign B[235] = \ML_int[9][235] ;
  assign B[234] = \ML_int[9][234] ;
  assign B[233] = \ML_int[9][233] ;
  assign B[232] = \ML_int[9][232] ;
  assign B[231] = \ML_int[9][231] ;
  assign B[230] = \ML_int[9][230] ;
  assign B[229] = \ML_int[9][229] ;
  assign B[228] = \ML_int[9][228] ;
  assign B[227] = \ML_int[9][227] ;
  assign B[226] = \ML_int[9][226] ;
  assign B[225] = \ML_int[9][225] ;
  assign B[224] = \ML_int[9][224] ;
  assign B[223] = \ML_int[9][223] ;
  assign B[222] = \ML_int[9][222] ;
  assign B[221] = \ML_int[9][221] ;
  assign B[220] = \ML_int[9][220] ;
  assign B[219] = \ML_int[9][219] ;
  assign B[218] = \ML_int[9][218] ;
  assign B[217] = \ML_int[9][217] ;
  assign B[216] = \ML_int[9][216] ;
  assign B[215] = \ML_int[9][215] ;
  assign B[214] = \ML_int[9][214] ;
  assign B[213] = \ML_int[9][213] ;
  assign B[212] = \ML_int[9][212] ;
  assign B[211] = \ML_int[9][211] ;
  assign B[210] = \ML_int[9][210] ;
  assign B[209] = \ML_int[9][209] ;
  assign B[208] = \ML_int[9][208] ;
  assign B[207] = \ML_int[9][207] ;
  assign B[206] = \ML_int[9][206] ;
  assign B[205] = \ML_int[9][205] ;
  assign B[204] = \ML_int[9][204] ;
  assign B[203] = \ML_int[9][203] ;
  assign B[202] = \ML_int[9][202] ;
  assign B[201] = \ML_int[9][201] ;
  assign B[200] = \ML_int[9][200] ;
  assign B[199] = \ML_int[9][199] ;
  assign B[198] = \ML_int[9][198] ;
  assign B[197] = \ML_int[9][197] ;
  assign B[196] = \ML_int[9][196] ;
  assign B[195] = \ML_int[9][195] ;
  assign B[194] = \ML_int[9][194] ;
  assign B[193] = \ML_int[9][193] ;
  assign B[192] = \ML_int[9][192] ;
  assign B[191] = \ML_int[9][191] ;
  assign B[190] = \ML_int[9][190] ;
  assign B[189] = \ML_int[9][189] ;
  assign B[188] = \ML_int[9][188] ;
  assign B[187] = \ML_int[9][187] ;
  assign B[186] = \ML_int[9][186] ;
  assign B[185] = \ML_int[9][185] ;
  assign B[184] = \ML_int[9][184] ;
  assign B[183] = \ML_int[9][183] ;
  assign B[182] = \ML_int[9][182] ;
  assign B[181] = \ML_int[9][181] ;
  assign B[180] = \ML_int[9][180] ;
  assign B[179] = \ML_int[9][179] ;
  assign B[178] = \ML_int[9][178] ;
  assign B[177] = \ML_int[9][177] ;
  assign B[176] = \ML_int[9][176] ;
  assign B[175] = \ML_int[9][175] ;
  assign B[174] = \ML_int[9][174] ;
  assign B[173] = \ML_int[9][173] ;
  assign B[172] = \ML_int[9][172] ;
  assign B[171] = \ML_int[9][171] ;
  assign B[170] = \ML_int[9][170] ;
  assign B[169] = \ML_int[9][169] ;
  assign B[168] = \ML_int[9][168] ;
  assign B[167] = \ML_int[9][167] ;
  assign B[166] = \ML_int[9][166] ;
  assign B[165] = \ML_int[9][165] ;
  assign B[164] = \ML_int[9][164] ;
  assign B[163] = \ML_int[9][163] ;
  assign B[162] = \ML_int[9][162] ;
  assign B[161] = \ML_int[9][161] ;
  assign B[160] = \ML_int[9][160] ;
  assign B[159] = \ML_int[9][159] ;
  assign B[158] = \ML_int[9][158] ;
  assign B[157] = \ML_int[9][157] ;
  assign B[156] = \ML_int[9][156] ;
  assign B[155] = \ML_int[9][155] ;
  assign B[154] = \ML_int[9][154] ;
  assign B[153] = \ML_int[9][153] ;
  assign B[152] = \ML_int[9][152] ;
  assign B[151] = \ML_int[9][151] ;
  assign B[150] = \ML_int[9][150] ;
  assign B[149] = \ML_int[9][149] ;
  assign B[148] = \ML_int[9][148] ;
  assign B[147] = \ML_int[9][147] ;
  assign B[146] = \ML_int[9][146] ;
  assign B[145] = \ML_int[9][145] ;
  assign B[144] = \ML_int[9][144] ;
  assign B[143] = \ML_int[9][143] ;
  assign B[142] = \ML_int[9][142] ;
  assign B[141] = \ML_int[9][141] ;
  assign B[140] = \ML_int[9][140] ;
  assign B[139] = \ML_int[9][139] ;
  assign B[138] = \ML_int[9][138] ;
  assign B[137] = \ML_int[9][137] ;
  assign B[136] = \ML_int[9][136] ;
  assign B[135] = \ML_int[9][135] ;
  assign B[134] = \ML_int[9][134] ;
  assign B[133] = \ML_int[9][133] ;
  assign B[132] = \ML_int[9][132] ;
  assign B[131] = \ML_int[9][131] ;
  assign B[130] = \ML_int[9][130] ;
  assign B[129] = \ML_int[9][129] ;
  assign B[128] = \ML_int[9][128] ;
  assign B[127] = \ML_int[9][127] ;
  assign B[126] = \ML_int[9][126] ;
  assign B[125] = \ML_int[9][125] ;
  assign B[124] = \ML_int[9][124] ;
  assign B[123] = \ML_int[9][123] ;
  assign B[122] = \ML_int[9][122] ;
  assign B[121] = \ML_int[9][121] ;
  assign B[120] = \ML_int[9][120] ;
  assign B[119] = \ML_int[9][119] ;
  assign B[118] = \ML_int[9][118] ;
  assign B[117] = \ML_int[9][117] ;
  assign B[116] = \ML_int[9][116] ;
  assign B[115] = \ML_int[9][115] ;
  assign B[114] = \ML_int[9][114] ;
  assign B[113] = \ML_int[9][113] ;
  assign B[112] = \ML_int[9][112] ;
  assign B[111] = \ML_int[9][111] ;
  assign B[110] = \ML_int[9][110] ;
  assign B[109] = \ML_int[9][109] ;
  assign B[108] = \ML_int[9][108] ;
  assign B[107] = \ML_int[9][107] ;
  assign B[106] = \ML_int[9][106] ;
  assign B[105] = \ML_int[9][105] ;
  assign B[104] = \ML_int[9][104] ;
  assign B[103] = \ML_int[9][103] ;
  assign B[102] = \ML_int[9][102] ;
  assign B[101] = \ML_int[9][101] ;
  assign B[100] = \ML_int[9][100] ;
  assign B[99] = \ML_int[9][99] ;
  assign B[98] = \ML_int[9][98] ;
  assign B[97] = \ML_int[9][97] ;
  assign B[96] = \ML_int[9][96] ;
  assign B[95] = \ML_int[9][95] ;
  assign B[94] = \ML_int[9][94] ;
  assign B[93] = \ML_int[9][93] ;
  assign B[92] = \ML_int[9][92] ;
  assign B[91] = \ML_int[9][91] ;
  assign B[90] = \ML_int[9][90] ;
  assign B[89] = \ML_int[9][89] ;
  assign B[88] = \ML_int[9][88] ;
  assign B[87] = \ML_int[9][87] ;
  assign B[86] = \ML_int[9][86] ;
  assign B[85] = \ML_int[9][85] ;
  assign B[84] = \ML_int[9][84] ;
  assign B[83] = \ML_int[9][83] ;
  assign B[82] = \ML_int[9][82] ;
  assign B[81] = \ML_int[9][81] ;
  assign B[80] = \ML_int[9][80] ;
  assign B[79] = \ML_int[9][79] ;
  assign B[78] = \ML_int[9][78] ;
  assign B[77] = \ML_int[9][77] ;
  assign B[76] = \ML_int[9][76] ;
  assign B[75] = \ML_int[9][75] ;
  assign B[74] = \ML_int[9][74] ;
  assign B[73] = \ML_int[9][73] ;
  assign B[72] = \ML_int[9][72] ;
  assign B[71] = \ML_int[9][71] ;
  assign B[70] = \ML_int[9][70] ;
  assign B[69] = \ML_int[9][69] ;
  assign B[68] = \ML_int[9][68] ;
  assign B[67] = \ML_int[9][67] ;
  assign B[66] = \ML_int[9][66] ;
  assign B[65] = \ML_int[9][65] ;
  assign B[64] = \ML_int[9][64] ;
  assign B[63] = \ML_int[9][63] ;
  assign B[62] = \ML_int[9][62] ;
  assign B[61] = \ML_int[9][61] ;
  assign B[60] = \ML_int[9][60] ;
  assign B[59] = \ML_int[9][59] ;
  assign B[58] = \ML_int[9][58] ;
  assign B[57] = \ML_int[9][57] ;
  assign B[56] = \ML_int[9][56] ;
  assign B[55] = \ML_int[9][55] ;
  assign B[54] = \ML_int[9][54] ;
  assign B[53] = \ML_int[9][53] ;
  assign B[52] = \ML_int[9][52] ;
  assign B[51] = \ML_int[9][51] ;
  assign B[50] = \ML_int[9][50] ;
  assign B[49] = \ML_int[9][49] ;
  assign B[48] = \ML_int[9][48] ;
  assign B[47] = \ML_int[9][47] ;
  assign B[46] = \ML_int[9][46] ;
  assign B[45] = \ML_int[9][45] ;
  assign B[44] = \ML_int[9][44] ;
  assign B[43] = \ML_int[9][43] ;
  assign B[42] = \ML_int[9][42] ;
  assign B[41] = \ML_int[9][41] ;
  assign B[40] = \ML_int[9][40] ;
  assign B[39] = \ML_int[9][39] ;
  assign B[38] = \ML_int[9][38] ;
  assign B[37] = \ML_int[9][37] ;
  assign B[36] = \ML_int[9][36] ;
  assign B[35] = \ML_int[9][35] ;
  assign B[34] = \ML_int[9][34] ;
  assign B[33] = \ML_int[9][33] ;
  assign B[32] = \ML_int[9][32] ;
  assign B[31] = \ML_int[9][31] ;
  assign B[30] = \ML_int[9][30] ;
  assign B[29] = \ML_int[9][29] ;
  assign B[28] = \ML_int[9][28] ;
  assign B[27] = \ML_int[9][27] ;
  assign B[26] = \ML_int[9][26] ;
  assign B[25] = \ML_int[9][25] ;
  assign B[24] = \ML_int[9][24] ;
  assign B[23] = \ML_int[9][23] ;
  assign B[22] = \ML_int[9][22] ;
  assign B[21] = \ML_int[9][21] ;
  assign B[20] = \ML_int[9][20] ;
  assign B[19] = \ML_int[9][19] ;
  assign B[18] = \ML_int[9][18] ;
  assign B[17] = \ML_int[9][17] ;
  assign B[16] = \ML_int[9][16] ;
  assign B[15] = \ML_int[9][15] ;
  assign B[14] = \ML_int[9][14] ;
  assign B[13] = \ML_int[9][13] ;
  assign B[12] = \ML_int[9][12] ;
  assign B[11] = \ML_int[9][11] ;
  assign B[10] = \ML_int[9][10] ;
  assign B[9] = \ML_int[9][9] ;
  assign B[8] = \ML_int[9][8] ;
  assign B[7] = \ML_int[9][7] ;
  assign B[6] = \ML_int[9][6] ;
  assign B[5] = \ML_int[9][5] ;
  assign B[4] = \ML_int[9][4] ;
  assign B[3] = \ML_int[9][3] ;
  assign B[2] = \ML_int[9][2] ;
  assign B[1] = \ML_int[9][1] ;
  assign B[0] = \ML_int[9][0] ;

  MUX2D1BWP M1_4_16 ( .I0(\MR_int[4][1] ), .I1(\ML_int[4][0] ), .S(SH[4]), .Z(
        \ML_int[5][16] ) );
  MUX2D1BWP M1_5_32 ( .I0(\ML_int[5][32] ), .I1(\ML_int[5][0] ), .S(SH[5]), 
        .Z(\ML_int[6][32] ) );
  MUX2D1BWP M1_6_64 ( .I0(\ML_int[6][64] ), .I1(\ML_int[6][0] ), .S(SH[6]), 
        .Z(\ML_int[7][64] ) );
  MUX2D1BWP M1_7_128 ( .I0(\ML_int[7][128] ), .I1(n26), .S(n21), .Z(
        \ML_int[8][128] ) );
  INVD1BWP U3 ( .I(n21), .ZN(n20) );
  INVD1BWP U4 ( .I(n22), .ZN(n19) );
  INVD1BWP U5 ( .I(n23), .ZN(n17) );
  INVD1BWP U6 ( .I(n22), .ZN(n18) );
  INVD1BWP U7 ( .I(n23), .ZN(n16) );
  INR2D1BWP U8 ( .A1(n33), .B1(n20), .ZN(\ML_int[8][177] ) );
  INVD1BWP U9 ( .I(n112), .ZN(n33) );
  INR2D1BWP U10 ( .A1(n29), .B1(n20), .ZN(\ML_int[8][176] ) );
  INVD1BWP U11 ( .I(n113), .ZN(n29) );
  INR2D1BWP U12 ( .A1(n31), .B1(n20), .ZN(\ML_int[8][161] ) );
  INVD1BWP U13 ( .I(n129), .ZN(n31) );
  INR2D1BWP U14 ( .A1(n27), .B1(n20), .ZN(\ML_int[8][160] ) );
  INVD1BWP U15 ( .I(n130), .ZN(n27) );
  INR2D1BWP U16 ( .A1(n32), .B1(n20), .ZN(\ML_int[8][145] ) );
  INVD1BWP U17 ( .I(n147), .ZN(n32) );
  INR2D1BWP U18 ( .A1(n28), .B1(n20), .ZN(\ML_int[8][144] ) );
  INVD1BWP U19 ( .I(n148), .ZN(n28) );
  INR2D1BWP U20 ( .A1(n34), .B1(n20), .ZN(\ML_int[8][130] ) );
  INVD1BWP U21 ( .I(n133), .ZN(n34) );
  INR2D1BWP U22 ( .A1(n30), .B1(n20), .ZN(\ML_int[8][129] ) );
  INVD1BWP U23 ( .I(n144), .ZN(n30) );
  INR2D1BWP U24 ( .A1(n87), .B1(n19), .ZN(\ML_int[8][191] ) );
  INVD1BWP U25 ( .I(n96), .ZN(n87) );
  INR2D1BWP U26 ( .A1(n73), .B1(n19), .ZN(\ML_int[8][190] ) );
  INVD1BWP U27 ( .I(n97), .ZN(n73) );
  INR2D1BWP U28 ( .A1(n77), .B1(n18), .ZN(\ML_int[8][189] ) );
  INVD1BWP U29 ( .I(n98), .ZN(n77) );
  INR2D1BWP U30 ( .A1(n81), .B1(n18), .ZN(\ML_int[8][188] ) );
  INVD1BWP U31 ( .I(n99), .ZN(n81) );
  INR2D1BWP U32 ( .A1(n85), .B1(n18), .ZN(\ML_int[8][187] ) );
  INVD1BWP U33 ( .I(n101), .ZN(n85) );
  INR2D1BWP U34 ( .A1(n69), .B1(n17), .ZN(\ML_int[8][186] ) );
  INVD1BWP U35 ( .I(n102), .ZN(n69) );
  INR2D1BWP U36 ( .A1(n65), .B1(n17), .ZN(\ML_int[8][185] ) );
  INVD1BWP U37 ( .I(n103), .ZN(n65) );
  INR2D1BWP U38 ( .A1(n61), .B1(n16), .ZN(\ML_int[8][184] ) );
  INVD1BWP U39 ( .I(n104), .ZN(n61) );
  INR2D1BWP U40 ( .A1(n57), .B1(n16), .ZN(\ML_int[8][183] ) );
  INVD1BWP U41 ( .I(n105), .ZN(n57) );
  INR2D1BWP U42 ( .A1(n53), .B1(n16), .ZN(\ML_int[8][182] ) );
  INVD1BWP U43 ( .I(n106), .ZN(n53) );
  INR2D1BWP U44 ( .A1(n49), .B1(n19), .ZN(\ML_int[8][181] ) );
  INVD1BWP U45 ( .I(n107), .ZN(n49) );
  INR2D1BWP U46 ( .A1(n45), .B1(n18), .ZN(\ML_int[8][180] ) );
  INVD1BWP U47 ( .I(n108), .ZN(n45) );
  INR2D1BWP U48 ( .A1(n89), .B1(n19), .ZN(\ML_int[8][175] ) );
  INVD1BWP U49 ( .I(n114), .ZN(n89) );
  INR2D1BWP U50 ( .A1(n71), .B1(n19), .ZN(\ML_int[8][174] ) );
  INVD1BWP U51 ( .I(n115), .ZN(n71) );
  INR2D1BWP U52 ( .A1(n75), .B1(n19), .ZN(\ML_int[8][173] ) );
  INVD1BWP U53 ( .I(n116), .ZN(n75) );
  INR2D1BWP U54 ( .A1(n79), .B1(n18), .ZN(\ML_int[8][172] ) );
  INVD1BWP U55 ( .I(n117), .ZN(n79) );
  INR2D1BWP U56 ( .A1(n83), .B1(n18), .ZN(\ML_int[8][171] ) );
  INVD1BWP U57 ( .I(n118), .ZN(n83) );
  INR2D1BWP U58 ( .A1(n67), .B1(n18), .ZN(\ML_int[8][170] ) );
  INVD1BWP U59 ( .I(n119), .ZN(n67) );
  INR2D1BWP U60 ( .A1(n63), .B1(n17), .ZN(\ML_int[8][169] ) );
  INVD1BWP U61 ( .I(n120), .ZN(n63) );
  INR2D1BWP U62 ( .A1(n59), .B1(n17), .ZN(\ML_int[8][168] ) );
  INVD1BWP U63 ( .I(n121), .ZN(n59) );
  INR2D1BWP U64 ( .A1(n55), .B1(n16), .ZN(\ML_int[8][167] ) );
  INVD1BWP U65 ( .I(n123), .ZN(n55) );
  INR2D1BWP U66 ( .A1(n51), .B1(n16), .ZN(\ML_int[8][166] ) );
  INVD1BWP U67 ( .I(n124), .ZN(n51) );
  INR2D1BWP U68 ( .A1(n47), .B1(n16), .ZN(\ML_int[8][165] ) );
  INVD1BWP U69 ( .I(n125), .ZN(n47) );
  INR2D1BWP U70 ( .A1(n43), .B1(n17), .ZN(\ML_int[8][164] ) );
  INVD1BWP U71 ( .I(n126), .ZN(n43) );
  INR2D1BWP U72 ( .A1(n86), .B1(n19), .ZN(\ML_int[8][159] ) );
  INVD1BWP U73 ( .I(n131), .ZN(n86) );
  INR2D1BWP U74 ( .A1(n72), .B1(n19), .ZN(\ML_int[8][158] ) );
  INVD1BWP U75 ( .I(n132), .ZN(n72) );
  INR2D1BWP U76 ( .A1(n76), .B1(n18), .ZN(\ML_int[8][157] ) );
  INVD1BWP U77 ( .I(n134), .ZN(n76) );
  INR2D1BWP U78 ( .A1(n80), .B1(n18), .ZN(\ML_int[8][156] ) );
  INVD1BWP U79 ( .I(n135), .ZN(n80) );
  INR2D1BWP U80 ( .A1(n84), .B1(n18), .ZN(\ML_int[8][155] ) );
  INVD1BWP U81 ( .I(n136), .ZN(n84) );
  INR2D1BWP U82 ( .A1(n68), .B1(n17), .ZN(\ML_int[8][154] ) );
  INVD1BWP U83 ( .I(n137), .ZN(n68) );
  INR2D1BWP U84 ( .A1(n64), .B1(n17), .ZN(\ML_int[8][153] ) );
  INVD1BWP U85 ( .I(n138), .ZN(n64) );
  INR2D1BWP U86 ( .A1(n60), .B1(n17), .ZN(\ML_int[8][152] ) );
  INVD1BWP U87 ( .I(n139), .ZN(n60) );
  INR2D1BWP U88 ( .A1(n56), .B1(n16), .ZN(\ML_int[8][151] ) );
  INVD1BWP U89 ( .I(n140), .ZN(n56) );
  INR2D1BWP U90 ( .A1(n52), .B1(n16), .ZN(\ML_int[8][150] ) );
  INVD1BWP U91 ( .I(n141), .ZN(n52) );
  INR2D1BWP U92 ( .A1(n48), .B1(n16), .ZN(\ML_int[8][149] ) );
  INVD1BWP U93 ( .I(n142), .ZN(n48) );
  INR2D1BWP U94 ( .A1(n44), .B1(n18), .ZN(\ML_int[8][148] ) );
  INVD1BWP U95 ( .I(n143), .ZN(n44) );
  INR2D1BWP U96 ( .A1(n88), .B1(n19), .ZN(\ML_int[8][143] ) );
  INVD1BWP U97 ( .I(n149), .ZN(n88) );
  INR2D1BWP U98 ( .A1(n70), .B1(n19), .ZN(\ML_int[8][142] ) );
  INVD1BWP U99 ( .I(n150), .ZN(n70) );
  INR2D1BWP U100 ( .A1(n74), .B1(n19), .ZN(\ML_int[8][141] ) );
  INVD1BWP U101 ( .I(n151), .ZN(n74) );
  INR2D1BWP U102 ( .A1(n78), .B1(n18), .ZN(\ML_int[8][140] ) );
  INVD1BWP U103 ( .I(n152), .ZN(n78) );
  INR2D1BWP U104 ( .A1(n82), .B1(n18), .ZN(\ML_int[8][139] ) );
  INVD1BWP U105 ( .I(n153), .ZN(n82) );
  INR2D1BWP U106 ( .A1(n66), .B1(n17), .ZN(\ML_int[8][138] ) );
  INVD1BWP U107 ( .I(n154), .ZN(n66) );
  INR2D1BWP U108 ( .A1(n62), .B1(n17), .ZN(\ML_int[8][137] ) );
  INVD1BWP U109 ( .I(n92), .ZN(n62) );
  INR2D1BWP U110 ( .A1(n58), .B1(n17), .ZN(\ML_int[8][136] ) );
  INVD1BWP U111 ( .I(n93), .ZN(n58) );
  INR2D1BWP U112 ( .A1(n54), .B1(n16), .ZN(\ML_int[8][135] ) );
  INVD1BWP U113 ( .I(n94), .ZN(n54) );
  INR2D1BWP U114 ( .A1(n50), .B1(n16), .ZN(\ML_int[8][134] ) );
  INVD1BWP U115 ( .I(n95), .ZN(n50) );
  INR2D1BWP U116 ( .A1(n46), .B1(n16), .ZN(\ML_int[8][133] ) );
  INVD1BWP U117 ( .I(n100), .ZN(n46) );
  INR2D1BWP U118 ( .A1(n42), .B1(n20), .ZN(\ML_int[8][132] ) );
  INVD1BWP U119 ( .I(n111), .ZN(n42) );
  INR2D1BWP U120 ( .A1(n41), .B1(n18), .ZN(\ML_int[8][179] ) );
  INVD1BWP U121 ( .I(n109), .ZN(n41) );
  INR2D1BWP U122 ( .A1(n37), .B1(n19), .ZN(\ML_int[8][178] ) );
  INVD1BWP U123 ( .I(n110), .ZN(n37) );
  INR2D1BWP U124 ( .A1(n39), .B1(n19), .ZN(\ML_int[8][163] ) );
  INVD1BWP U125 ( .I(n127), .ZN(n39) );
  INR2D1BWP U126 ( .A1(n35), .B1(n18), .ZN(\ML_int[8][162] ) );
  INVD1BWP U127 ( .I(n128), .ZN(n35) );
  INR2D1BWP U128 ( .A1(n40), .B1(n17), .ZN(\ML_int[8][147] ) );
  INVD1BWP U129 ( .I(n145), .ZN(n40) );
  INR2D1BWP U130 ( .A1(n36), .B1(n16), .ZN(\ML_int[8][146] ) );
  INVD1BWP U131 ( .I(n146), .ZN(n36) );
  INR2D1BWP U132 ( .A1(n38), .B1(n20), .ZN(\ML_int[8][131] ) );
  INVD1BWP U133 ( .I(n122), .ZN(n38) );
  CKBD1BWP U134 ( .I(n13), .Z(n6) );
  CKBD1BWP U135 ( .I(n13), .Z(n7) );
  CKBD1BWP U136 ( .I(n12), .Z(n10) );
  CKBD1BWP U137 ( .I(n12), .Z(n9) );
  CKBD1BWP U138 ( .I(n13), .Z(n8) );
  CKBD1BWP U139 ( .I(n14), .Z(n3) );
  CKBD1BWP U140 ( .I(n14), .Z(n4) );
  CKBD1BWP U141 ( .I(n14), .Z(n5) );
  CKBD1BWP U142 ( .I(n15), .Z(n1) );
  CKBD1BWP U143 ( .I(n15), .Z(n2) );
  CKBD1BWP U144 ( .I(n12), .Z(n11) );
  CKBD1BWP U145 ( .I(n91), .Z(n12) );
  CKBD1BWP U146 ( .I(n91), .Z(n13) );
  CKBD1BWP U147 ( .I(n91), .Z(n14) );
  CKBD1BWP U148 ( .I(n91), .Z(n15) );
  NR2XD0BWP U149 ( .A1(n24), .A2(n25), .ZN(\ML_int[7][128] ) );
  INVD1BWP U150 ( .I(n155), .ZN(n26) );
  INVD1BWP U151 ( .I(\ML_int[6][64] ), .ZN(n24) );
  INR2D1BWP U152 ( .A1(\ML_int[7][81] ), .B1(n20), .ZN(\ML_int[8][209] ) );
  INR2D1BWP U153 ( .A1(\ML_int[7][80] ), .B1(n20), .ZN(\ML_int[8][208] ) );
  INR2D1BWP U154 ( .A1(\ML_int[7][66] ), .B1(n20), .ZN(\ML_int[8][194] ) );
  INR2D1BWP U155 ( .A1(\ML_int[7][65] ), .B1(n20), .ZN(\ML_int[8][193] ) );
  INR2D1BWP U156 ( .A1(\ML_int[7][64] ), .B1(n20), .ZN(\ML_int[8][192] ) );
  INR2D1BWP U157 ( .A1(\ML_int[7][127] ), .B1(n20), .ZN(\ML_int[8][255] ) );
  INR2D1BWP U158 ( .A1(\ML_int[7][126] ), .B1(n16), .ZN(\ML_int[8][254] ) );
  INR2D1BWP U159 ( .A1(\ML_int[7][125] ), .B1(n19), .ZN(\ML_int[8][253] ) );
  INR2D1BWP U160 ( .A1(\ML_int[7][124] ), .B1(n18), .ZN(\ML_int[8][252] ) );
  INR2D1BWP U161 ( .A1(\ML_int[7][123] ), .B1(n17), .ZN(\ML_int[8][251] ) );
  INR2D1BWP U162 ( .A1(\ML_int[7][122] ), .B1(n19), .ZN(\ML_int[8][250] ) );
  INR2D1BWP U163 ( .A1(\ML_int[7][121] ), .B1(n20), .ZN(\ML_int[8][249] ) );
  INR2D1BWP U164 ( .A1(\ML_int[7][120] ), .B1(n18), .ZN(\ML_int[8][248] ) );
  INR2D1BWP U165 ( .A1(\ML_int[7][119] ), .B1(n17), .ZN(\ML_int[8][247] ) );
  INR2D1BWP U166 ( .A1(\ML_int[7][118] ), .B1(n16), .ZN(\ML_int[8][246] ) );
  INR2D1BWP U167 ( .A1(\ML_int[7][117] ), .B1(n19), .ZN(\ML_int[8][245] ) );
  INR2D1BWP U168 ( .A1(\ML_int[7][116] ), .B1(n20), .ZN(\ML_int[8][244] ) );
  INR2D1BWP U169 ( .A1(\ML_int[7][115] ), .B1(n18), .ZN(\ML_int[8][243] ) );
  INR2D1BWP U170 ( .A1(\ML_int[7][114] ), .B1(n17), .ZN(\ML_int[8][242] ) );
  INR2D1BWP U171 ( .A1(\ML_int[7][113] ), .B1(n16), .ZN(\ML_int[8][241] ) );
  INR2D1BWP U172 ( .A1(\ML_int[7][112] ), .B1(n19), .ZN(\ML_int[8][240] ) );
  INR2D1BWP U173 ( .A1(\ML_int[7][111] ), .B1(n20), .ZN(\ML_int[8][239] ) );
  INR2D1BWP U174 ( .A1(\ML_int[7][110] ), .B1(n18), .ZN(\ML_int[8][238] ) );
  INR2D1BWP U175 ( .A1(\ML_int[7][109] ), .B1(n20), .ZN(\ML_int[8][237] ) );
  INR2D1BWP U176 ( .A1(\ML_int[7][108] ), .B1(n18), .ZN(\ML_int[8][236] ) );
  INR2D1BWP U177 ( .A1(\ML_int[7][107] ), .B1(n17), .ZN(\ML_int[8][235] ) );
  INR2D1BWP U178 ( .A1(\ML_int[7][106] ), .B1(n16), .ZN(\ML_int[8][234] ) );
  INR2D1BWP U179 ( .A1(\ML_int[7][105] ), .B1(n17), .ZN(\ML_int[8][233] ) );
  INR2D1BWP U180 ( .A1(\ML_int[7][104] ), .B1(n19), .ZN(\ML_int[8][232] ) );
  INR2D1BWP U181 ( .A1(\ML_int[7][103] ), .B1(n20), .ZN(\ML_int[8][231] ) );
  INR2D1BWP U182 ( .A1(\ML_int[7][102] ), .B1(n18), .ZN(\ML_int[8][230] ) );
  INR2D1BWP U183 ( .A1(\ML_int[7][101] ), .B1(n17), .ZN(\ML_int[8][229] ) );
  INR2D1BWP U184 ( .A1(\ML_int[7][100] ), .B1(n16), .ZN(\ML_int[8][228] ) );
  INR2D1BWP U185 ( .A1(\ML_int[7][99] ), .B1(n16), .ZN(\ML_int[8][227] ) );
  INR2D1BWP U186 ( .A1(\ML_int[7][98] ), .B1(n19), .ZN(\ML_int[8][226] ) );
  INR2D1BWP U187 ( .A1(\ML_int[7][97] ), .B1(n20), .ZN(\ML_int[8][225] ) );
  INR2D1BWP U188 ( .A1(\ML_int[7][96] ), .B1(n18), .ZN(\ML_int[8][224] ) );
  INR2D1BWP U189 ( .A1(\ML_int[7][95] ), .B1(n17), .ZN(\ML_int[8][223] ) );
  INR2D1BWP U190 ( .A1(\ML_int[7][94] ), .B1(n16), .ZN(\ML_int[8][222] ) );
  INR2D1BWP U191 ( .A1(\ML_int[7][93] ), .B1(n19), .ZN(\ML_int[8][221] ) );
  INR2D1BWP U192 ( .A1(\ML_int[7][92] ), .B1(n18), .ZN(\ML_int[8][220] ) );
  INR2D1BWP U193 ( .A1(\ML_int[7][91] ), .B1(n20), .ZN(\ML_int[8][219] ) );
  INR2D1BWP U194 ( .A1(\ML_int[7][90] ), .B1(n19), .ZN(\ML_int[8][218] ) );
  INR2D1BWP U195 ( .A1(\ML_int[7][89] ), .B1(n18), .ZN(\ML_int[8][217] ) );
  INR2D1BWP U196 ( .A1(\ML_int[7][88] ), .B1(n17), .ZN(\ML_int[8][216] ) );
  INR2D1BWP U197 ( .A1(\ML_int[7][87] ), .B1(n16), .ZN(\ML_int[8][215] ) );
  INR2D1BWP U198 ( .A1(\ML_int[7][86] ), .B1(n20), .ZN(\ML_int[8][214] ) );
  INR2D1BWP U199 ( .A1(\ML_int[7][85] ), .B1(n17), .ZN(\ML_int[8][213] ) );
  INR2D1BWP U200 ( .A1(\ML_int[7][84] ), .B1(n20), .ZN(\ML_int[8][212] ) );
  INR2D1BWP U201 ( .A1(\ML_int[7][79] ), .B1(n19), .ZN(\ML_int[8][207] ) );
  INR2D1BWP U202 ( .A1(\ML_int[7][78] ), .B1(n19), .ZN(\ML_int[8][206] ) );
  INR2D1BWP U203 ( .A1(\ML_int[7][77] ), .B1(n19), .ZN(\ML_int[8][205] ) );
  INR2D1BWP U204 ( .A1(\ML_int[7][76] ), .B1(n18), .ZN(\ML_int[8][204] ) );
  INR2D1BWP U205 ( .A1(\ML_int[7][75] ), .B1(n18), .ZN(\ML_int[8][203] ) );
  INR2D1BWP U206 ( .A1(\ML_int[7][74] ), .B1(n17), .ZN(\ML_int[8][202] ) );
  INR2D1BWP U207 ( .A1(\ML_int[7][73] ), .B1(n17), .ZN(\ML_int[8][201] ) );
  INR2D1BWP U208 ( .A1(\ML_int[7][72] ), .B1(n17), .ZN(\ML_int[8][200] ) );
  INR2D1BWP U209 ( .A1(\ML_int[7][71] ), .B1(n16), .ZN(\ML_int[8][199] ) );
  INR2D1BWP U210 ( .A1(\ML_int[7][70] ), .B1(n16), .ZN(\ML_int[8][198] ) );
  INR2D1BWP U211 ( .A1(\ML_int[7][69] ), .B1(n16), .ZN(\ML_int[8][197] ) );
  INR2D1BWP U212 ( .A1(\ML_int[7][68] ), .B1(n17), .ZN(\ML_int[8][196] ) );
  INR2D1BWP U213 ( .A1(\ML_int[7][83] ), .B1(n16), .ZN(\ML_int[8][211] ) );
  INR2D1BWP U214 ( .A1(\ML_int[7][82] ), .B1(n20), .ZN(\ML_int[8][210] ) );
  INR2D1BWP U215 ( .A1(\ML_int[7][67] ), .B1(n19), .ZN(\ML_int[8][195] ) );
  INVD1BWP U216 ( .I(SH[6]), .ZN(n90) );
  INVD1BWP U217 ( .I(SH[6]), .ZN(n25) );
  AN2XD1BWP U218 ( .A1(\ML_int[6][63] ), .A2(SH[6]), .Z(\ML_int[7][127] ) );
  AN2XD1BWP U219 ( .A1(\ML_int[6][62] ), .A2(SH[6]), .Z(\ML_int[7][126] ) );
  AN2XD1BWP U220 ( .A1(\ML_int[6][61] ), .A2(SH[6]), .Z(\ML_int[7][125] ) );
  AN2XD1BWP U221 ( .A1(\ML_int[6][60] ), .A2(SH[6]), .Z(\ML_int[7][124] ) );
  AN2XD1BWP U222 ( .A1(\ML_int[6][59] ), .A2(SH[6]), .Z(\ML_int[7][123] ) );
  AN2XD1BWP U223 ( .A1(\ML_int[6][58] ), .A2(SH[6]), .Z(\ML_int[7][122] ) );
  AN2XD1BWP U224 ( .A1(\ML_int[6][57] ), .A2(SH[6]), .Z(\ML_int[7][121] ) );
  AN2XD1BWP U225 ( .A1(\ML_int[6][56] ), .A2(SH[6]), .Z(\ML_int[7][120] ) );
  AN2XD1BWP U226 ( .A1(\ML_int[6][55] ), .A2(SH[6]), .Z(\ML_int[7][119] ) );
  AN2XD1BWP U227 ( .A1(\ML_int[6][54] ), .A2(SH[6]), .Z(\ML_int[7][118] ) );
  AN2XD1BWP U228 ( .A1(\ML_int[6][53] ), .A2(SH[6]), .Z(\ML_int[7][117] ) );
  AN2XD1BWP U229 ( .A1(\ML_int[6][52] ), .A2(SH[6]), .Z(\ML_int[7][116] ) );
  AN2XD1BWP U230 ( .A1(\ML_int[6][51] ), .A2(SH[6]), .Z(\ML_int[7][115] ) );
  AN2XD1BWP U231 ( .A1(\ML_int[6][50] ), .A2(SH[6]), .Z(\ML_int[7][114] ) );
  AN2XD1BWP U232 ( .A1(\ML_int[6][49] ), .A2(SH[6]), .Z(\ML_int[7][113] ) );
  AN2XD1BWP U233 ( .A1(\ML_int[6][48] ), .A2(SH[6]), .Z(\ML_int[7][112] ) );
  AN2XD1BWP U234 ( .A1(\ML_int[6][47] ), .A2(SH[6]), .Z(\ML_int[7][111] ) );
  AN2XD1BWP U235 ( .A1(\ML_int[6][46] ), .A2(SH[6]), .Z(\ML_int[7][110] ) );
  AN2XD1BWP U236 ( .A1(\ML_int[6][45] ), .A2(SH[6]), .Z(\ML_int[7][109] ) );
  AN2XD1BWP U237 ( .A1(\ML_int[6][44] ), .A2(SH[6]), .Z(\ML_int[7][108] ) );
  AN2XD1BWP U238 ( .A1(\ML_int[6][43] ), .A2(SH[6]), .Z(\ML_int[7][107] ) );
  AN2XD1BWP U239 ( .A1(\ML_int[6][42] ), .A2(SH[6]), .Z(\ML_int[7][106] ) );
  AN2XD1BWP U240 ( .A1(\ML_int[6][41] ), .A2(SH[6]), .Z(\ML_int[7][105] ) );
  AN2XD1BWP U241 ( .A1(\ML_int[6][40] ), .A2(SH[6]), .Z(\ML_int[7][104] ) );
  AN2XD1BWP U242 ( .A1(\ML_int[6][39] ), .A2(SH[6]), .Z(\ML_int[7][103] ) );
  AN2XD1BWP U243 ( .A1(\ML_int[6][38] ), .A2(SH[6]), .Z(\ML_int[7][102] ) );
  AN2XD1BWP U244 ( .A1(\ML_int[6][37] ), .A2(SH[6]), .Z(\ML_int[7][101] ) );
  AN2XD1BWP U245 ( .A1(\ML_int[6][36] ), .A2(SH[6]), .Z(\ML_int[7][100] ) );
  AN2XD1BWP U246 ( .A1(\ML_int[6][35] ), .A2(SH[6]), .Z(\ML_int[7][99] ) );
  AN2XD1BWP U247 ( .A1(\ML_int[6][34] ), .A2(SH[6]), .Z(\ML_int[7][98] ) );
  AN2XD1BWP U248 ( .A1(\ML_int[6][33] ), .A2(SH[6]), .Z(\ML_int[7][97] ) );
  AN2XD1BWP U249 ( .A1(\ML_int[6][32] ), .A2(SH[6]), .Z(\ML_int[7][96] ) );
  AN2XD1BWP U250 ( .A1(\ML_int[6][31] ), .A2(SH[6]), .Z(\ML_int[7][95] ) );
  AN2XD1BWP U251 ( .A1(\ML_int[6][30] ), .A2(SH[6]), .Z(\ML_int[7][94] ) );
  AN2XD1BWP U252 ( .A1(\ML_int[6][29] ), .A2(SH[6]), .Z(\ML_int[7][93] ) );
  AN2XD1BWP U253 ( .A1(\ML_int[6][28] ), .A2(SH[6]), .Z(\ML_int[7][92] ) );
  AN2XD1BWP U254 ( .A1(\ML_int[6][27] ), .A2(SH[6]), .Z(\ML_int[7][91] ) );
  AN2XD1BWP U255 ( .A1(\ML_int[6][26] ), .A2(SH[6]), .Z(\ML_int[7][90] ) );
  AN2XD1BWP U256 ( .A1(\ML_int[6][25] ), .A2(SH[6]), .Z(\ML_int[7][89] ) );
  AN2XD1BWP U257 ( .A1(\ML_int[6][24] ), .A2(SH[6]), .Z(\ML_int[7][88] ) );
  AN2XD1BWP U258 ( .A1(\ML_int[6][23] ), .A2(SH[6]), .Z(\ML_int[7][87] ) );
  AN2XD1BWP U259 ( .A1(\ML_int[6][22] ), .A2(SH[6]), .Z(\ML_int[7][86] ) );
  AN2XD1BWP U260 ( .A1(\ML_int[6][21] ), .A2(SH[6]), .Z(\ML_int[7][85] ) );
  AN2XD1BWP U261 ( .A1(\ML_int[6][20] ), .A2(SH[6]), .Z(\ML_int[7][84] ) );
  AN2XD1BWP U262 ( .A1(\ML_int[6][19] ), .A2(SH[6]), .Z(\ML_int[7][83] ) );
  AN2XD1BWP U263 ( .A1(\ML_int[6][18] ), .A2(SH[6]), .Z(\ML_int[7][82] ) );
  AN2XD1BWP U264 ( .A1(\ML_int[6][17] ), .A2(SH[6]), .Z(\ML_int[7][81] ) );
  AN2XD1BWP U265 ( .A1(\ML_int[6][16] ), .A2(SH[6]), .Z(\ML_int[7][80] ) );
  AN2XD1BWP U266 ( .A1(\ML_int[6][15] ), .A2(SH[6]), .Z(\ML_int[7][79] ) );
  AN2XD1BWP U267 ( .A1(\ML_int[6][14] ), .A2(SH[6]), .Z(\ML_int[7][78] ) );
  AN2XD1BWP U268 ( .A1(\ML_int[6][13] ), .A2(SH[6]), .Z(\ML_int[7][77] ) );
  AN2XD1BWP U269 ( .A1(\ML_int[6][12] ), .A2(SH[6]), .Z(\ML_int[7][76] ) );
  AN2XD1BWP U270 ( .A1(\ML_int[6][11] ), .A2(SH[6]), .Z(\ML_int[7][75] ) );
  AN2XD1BWP U271 ( .A1(\ML_int[6][10] ), .A2(SH[6]), .Z(\ML_int[7][74] ) );
  AN2XD1BWP U272 ( .A1(\ML_int[6][9] ), .A2(SH[6]), .Z(\ML_int[7][73] ) );
  AN2XD1BWP U273 ( .A1(\ML_int[6][8] ), .A2(SH[6]), .Z(\ML_int[7][72] ) );
  AN2XD1BWP U274 ( .A1(\ML_int[6][7] ), .A2(SH[6]), .Z(\ML_int[7][71] ) );
  AN2XD1BWP U275 ( .A1(\ML_int[6][6] ), .A2(SH[6]), .Z(\ML_int[7][70] ) );
  AN2XD1BWP U276 ( .A1(\ML_int[6][5] ), .A2(SH[6]), .Z(\ML_int[7][69] ) );
  AN2XD1BWP U277 ( .A1(\ML_int[6][4] ), .A2(SH[6]), .Z(\ML_int[7][68] ) );
  AN2XD1BWP U278 ( .A1(\ML_int[6][3] ), .A2(SH[6]), .Z(\ML_int[7][67] ) );
  AN2XD1BWP U279 ( .A1(\ML_int[6][2] ), .A2(SH[6]), .Z(\ML_int[7][66] ) );
  AN2XD1BWP U280 ( .A1(\ML_int[6][1] ), .A2(SH[6]), .Z(\ML_int[7][65] ) );
  AN2XD1BWP U281 ( .A1(\ML_int[5][32] ), .A2(SH[5]), .Z(\ML_int[6][64] ) );
  AN2XD1BWP U282 ( .A1(\ML_int[5][31] ), .A2(SH[5]), .Z(\ML_int[6][63] ) );
  AN2XD1BWP U283 ( .A1(\ML_int[5][30] ), .A2(SH[5]), .Z(\ML_int[6][62] ) );
  AN2XD1BWP U284 ( .A1(\ML_int[5][29] ), .A2(SH[5]), .Z(\ML_int[6][61] ) );
  AN2XD1BWP U285 ( .A1(\ML_int[5][28] ), .A2(SH[5]), .Z(\ML_int[6][60] ) );
  AN2XD1BWP U286 ( .A1(\ML_int[5][27] ), .A2(SH[5]), .Z(\ML_int[6][59] ) );
  AN2XD1BWP U287 ( .A1(\ML_int[5][26] ), .A2(SH[5]), .Z(\ML_int[6][58] ) );
  AN2XD1BWP U288 ( .A1(\ML_int[5][25] ), .A2(SH[5]), .Z(\ML_int[6][57] ) );
  AN2XD1BWP U289 ( .A1(\ML_int[5][24] ), .A2(SH[5]), .Z(\ML_int[6][56] ) );
  AN2XD1BWP U290 ( .A1(\ML_int[5][23] ), .A2(SH[5]), .Z(\ML_int[6][55] ) );
  AN2XD1BWP U291 ( .A1(\ML_int[5][22] ), .A2(SH[5]), .Z(\ML_int[6][54] ) );
  AN2XD1BWP U292 ( .A1(\ML_int[5][21] ), .A2(SH[5]), .Z(\ML_int[6][53] ) );
  AN2XD1BWP U293 ( .A1(\ML_int[5][20] ), .A2(SH[5]), .Z(\ML_int[6][52] ) );
  AN2XD1BWP U294 ( .A1(\ML_int[5][19] ), .A2(SH[5]), .Z(\ML_int[6][51] ) );
  AN2XD1BWP U295 ( .A1(\ML_int[5][18] ), .A2(SH[5]), .Z(\ML_int[6][50] ) );
  AN2XD1BWP U296 ( .A1(\ML_int[5][17] ), .A2(SH[5]), .Z(\ML_int[6][49] ) );
  AN2XD1BWP U297 ( .A1(\ML_int[5][16] ), .A2(SH[5]), .Z(\ML_int[6][48] ) );
  AN2XD1BWP U298 ( .A1(\ML_int[5][15] ), .A2(SH[5]), .Z(\ML_int[6][47] ) );
  AN2XD1BWP U299 ( .A1(\ML_int[5][14] ), .A2(SH[5]), .Z(\ML_int[6][46] ) );
  AN2XD1BWP U300 ( .A1(\ML_int[5][13] ), .A2(SH[5]), .Z(\ML_int[6][45] ) );
  AN2XD1BWP U301 ( .A1(\ML_int[5][12] ), .A2(SH[5]), .Z(\ML_int[6][44] ) );
  AN2XD1BWP U302 ( .A1(\ML_int[5][11] ), .A2(SH[5]), .Z(\ML_int[6][43] ) );
  AN2XD1BWP U303 ( .A1(\ML_int[5][10] ), .A2(SH[5]), .Z(\ML_int[6][42] ) );
  AN2XD1BWP U304 ( .A1(\ML_int[5][9] ), .A2(SH[5]), .Z(\ML_int[6][41] ) );
  AN2XD1BWP U305 ( .A1(\ML_int[5][8] ), .A2(SH[5]), .Z(\ML_int[6][40] ) );
  AN2XD1BWP U306 ( .A1(\ML_int[5][7] ), .A2(SH[5]), .Z(\ML_int[6][39] ) );
  AN2XD1BWP U307 ( .A1(\ML_int[5][6] ), .A2(SH[5]), .Z(\ML_int[6][38] ) );
  AN2XD1BWP U308 ( .A1(\ML_int[5][5] ), .A2(SH[5]), .Z(\ML_int[6][37] ) );
  AN2XD1BWP U309 ( .A1(\ML_int[5][4] ), .A2(SH[5]), .Z(\ML_int[6][36] ) );
  AN2XD1BWP U310 ( .A1(\ML_int[5][3] ), .A2(SH[5]), .Z(\ML_int[6][35] ) );
  AN2XD1BWP U311 ( .A1(\ML_int[5][2] ), .A2(SH[5]), .Z(\ML_int[6][34] ) );
  AN2XD1BWP U312 ( .A1(\ML_int[5][1] ), .A2(SH[5]), .Z(\ML_int[6][33] ) );
  AN2XD1BWP U313 ( .A1(\MR_int[4][1] ), .A2(SH[4]), .Z(\ML_int[5][32] ) );
  AN2XD1BWP U314 ( .A1(\MR_int[4][0] ), .A2(SH[4]), .Z(\ML_int[5][31] ) );
  AN2XD1BWP U315 ( .A1(\ML_int[4][14] ), .A2(SH[4]), .Z(\ML_int[5][30] ) );
  AN2XD1BWP U316 ( .A1(\ML_int[4][13] ), .A2(SH[4]), .Z(\ML_int[5][29] ) );
  AN2XD1BWP U317 ( .A1(\ML_int[4][12] ), .A2(SH[4]), .Z(\ML_int[5][28] ) );
  AN2XD1BWP U318 ( .A1(\ML_int[4][11] ), .A2(SH[4]), .Z(\ML_int[5][27] ) );
  AN2XD1BWP U319 ( .A1(\ML_int[4][10] ), .A2(SH[4]), .Z(\ML_int[5][26] ) );
  AN2XD1BWP U320 ( .A1(\ML_int[4][9] ), .A2(SH[4]), .Z(\ML_int[5][25] ) );
  AN2XD1BWP U321 ( .A1(\ML_int[4][8] ), .A2(SH[4]), .Z(\ML_int[5][24] ) );
  AN2XD1BWP U322 ( .A1(\ML_int[4][7] ), .A2(SH[4]), .Z(\ML_int[5][23] ) );
  AN2XD1BWP U323 ( .A1(\ML_int[4][6] ), .A2(SH[4]), .Z(\ML_int[5][22] ) );
  AN2XD1BWP U324 ( .A1(\ML_int[4][5] ), .A2(SH[4]), .Z(\ML_int[5][21] ) );
  AN2XD1BWP U325 ( .A1(\ML_int[4][4] ), .A2(SH[4]), .Z(\ML_int[5][20] ) );
  AN2XD1BWP U326 ( .A1(\ML_int[4][3] ), .A2(SH[4]), .Z(\ML_int[5][19] ) );
  AN2XD1BWP U327 ( .A1(\ML_int[4][2] ), .A2(SH[4]), .Z(\ML_int[5][18] ) );
  AN2XD1BWP U328 ( .A1(\ML_int[4][1] ), .A2(SH[4]), .Z(\ML_int[5][17] ) );
  CKBD1BWP U329 ( .I(SH[7]), .Z(n21) );
  CKBD1BWP U330 ( .I(SH[7]), .Z(n22) );
  CKBD1BWP U331 ( .I(SH[7]), .Z(n23) );
  NR2D0BWP U332 ( .A1(n1), .A2(n92), .ZN(\ML_int[9][9] ) );
  INR2D0BWP U333 ( .A1(\ML_int[7][99] ), .B1(n11), .ZN(\ML_int[9][99] ) );
  INR2D0BWP U334 ( .A1(\ML_int[7][98] ), .B1(n11), .ZN(\ML_int[9][98] ) );
  INR2D0BWP U335 ( .A1(\ML_int[7][97] ), .B1(n10), .ZN(\ML_int[9][97] ) );
  INR2D0BWP U336 ( .A1(\ML_int[7][96] ), .B1(n10), .ZN(\ML_int[9][96] ) );
  INR2D0BWP U337 ( .A1(\ML_int[7][95] ), .B1(n10), .ZN(\ML_int[9][95] ) );
  INR2D0BWP U338 ( .A1(\ML_int[7][94] ), .B1(n10), .ZN(\ML_int[9][94] ) );
  INR2D0BWP U339 ( .A1(\ML_int[7][93] ), .B1(n10), .ZN(\ML_int[9][93] ) );
  INR2D0BWP U340 ( .A1(\ML_int[7][92] ), .B1(n10), .ZN(\ML_int[9][92] ) );
  INR2D0BWP U341 ( .A1(\ML_int[7][91] ), .B1(n10), .ZN(\ML_int[9][91] ) );
  INR2D0BWP U342 ( .A1(\ML_int[7][90] ), .B1(n10), .ZN(\ML_int[9][90] ) );
  NR2D0BWP U343 ( .A1(n1), .A2(n93), .ZN(\ML_int[9][8] ) );
  INR2D0BWP U344 ( .A1(\ML_int[7][89] ), .B1(n10), .ZN(\ML_int[9][89] ) );
  INR2D0BWP U345 ( .A1(\ML_int[7][88] ), .B1(n10), .ZN(\ML_int[9][88] ) );
  INR2D0BWP U346 ( .A1(\ML_int[7][87] ), .B1(n10), .ZN(\ML_int[9][87] ) );
  INR2D0BWP U347 ( .A1(\ML_int[7][86] ), .B1(n10), .ZN(\ML_int[9][86] ) );
  INR2D0BWP U348 ( .A1(\ML_int[7][85] ), .B1(n9), .ZN(\ML_int[9][85] ) );
  INR2D0BWP U349 ( .A1(\ML_int[7][84] ), .B1(n9), .ZN(\ML_int[9][84] ) );
  INR2D0BWP U350 ( .A1(\ML_int[7][83] ), .B1(n9), .ZN(\ML_int[9][83] ) );
  INR2D0BWP U351 ( .A1(\ML_int[7][82] ), .B1(n9), .ZN(\ML_int[9][82] ) );
  INR2D0BWP U352 ( .A1(\ML_int[7][81] ), .B1(n9), .ZN(\ML_int[9][81] ) );
  INR2D0BWP U353 ( .A1(\ML_int[7][80] ), .B1(n9), .ZN(\ML_int[9][80] ) );
  NR2D0BWP U354 ( .A1(n1), .A2(n94), .ZN(\ML_int[9][7] ) );
  INR2D0BWP U355 ( .A1(\ML_int[7][79] ), .B1(n9), .ZN(\ML_int[9][79] ) );
  INR2D0BWP U356 ( .A1(\ML_int[7][78] ), .B1(n9), .ZN(\ML_int[9][78] ) );
  INR2D0BWP U357 ( .A1(\ML_int[7][77] ), .B1(n9), .ZN(\ML_int[9][77] ) );
  INR2D0BWP U358 ( .A1(\ML_int[7][76] ), .B1(n9), .ZN(\ML_int[9][76] ) );
  INR2D0BWP U359 ( .A1(\ML_int[7][75] ), .B1(n9), .ZN(\ML_int[9][75] ) );
  INR2D0BWP U360 ( .A1(\ML_int[7][74] ), .B1(n9), .ZN(\ML_int[9][74] ) );
  INR2D0BWP U361 ( .A1(\ML_int[7][73] ), .B1(n8), .ZN(\ML_int[9][73] ) );
  INR2D0BWP U362 ( .A1(\ML_int[7][72] ), .B1(n8), .ZN(\ML_int[9][72] ) );
  INR2D0BWP U363 ( .A1(\ML_int[7][71] ), .B1(n8), .ZN(\ML_int[9][71] ) );
  INR2D0BWP U364 ( .A1(\ML_int[7][70] ), .B1(n8), .ZN(\ML_int[9][70] ) );
  NR2D0BWP U365 ( .A1(n1), .A2(n95), .ZN(\ML_int[9][6] ) );
  INR2D0BWP U366 ( .A1(\ML_int[7][69] ), .B1(n8), .ZN(\ML_int[9][69] ) );
  INR2D0BWP U367 ( .A1(\ML_int[7][68] ), .B1(n8), .ZN(\ML_int[9][68] ) );
  INR2D0BWP U368 ( .A1(\ML_int[7][67] ), .B1(n8), .ZN(\ML_int[9][67] ) );
  INR2D0BWP U369 ( .A1(\ML_int[7][66] ), .B1(n8), .ZN(\ML_int[9][66] ) );
  INR2D0BWP U370 ( .A1(\ML_int[7][65] ), .B1(n8), .ZN(\ML_int[9][65] ) );
  INR2D0BWP U371 ( .A1(\ML_int[7][64] ), .B1(n8), .ZN(\ML_int[9][64] ) );
  NR2D0BWP U372 ( .A1(n1), .A2(n96), .ZN(\ML_int[9][63] ) );
  NR2D0BWP U373 ( .A1(n1), .A2(n97), .ZN(\ML_int[9][62] ) );
  NR2D0BWP U374 ( .A1(n1), .A2(n98), .ZN(\ML_int[9][61] ) );
  NR2D0BWP U375 ( .A1(n1), .A2(n99), .ZN(\ML_int[9][60] ) );
  NR2D0BWP U376 ( .A1(n1), .A2(n100), .ZN(\ML_int[9][5] ) );
  NR2D0BWP U377 ( .A1(n1), .A2(n101), .ZN(\ML_int[9][59] ) );
  NR2D0BWP U378 ( .A1(n1), .A2(n102), .ZN(\ML_int[9][58] ) );
  NR2D0BWP U379 ( .A1(n1), .A2(n103), .ZN(\ML_int[9][57] ) );
  NR2D0BWP U380 ( .A1(n2), .A2(n104), .ZN(\ML_int[9][56] ) );
  NR2D0BWP U381 ( .A1(n2), .A2(n105), .ZN(\ML_int[9][55] ) );
  NR2D0BWP U382 ( .A1(n2), .A2(n106), .ZN(\ML_int[9][54] ) );
  NR2D0BWP U383 ( .A1(n2), .A2(n107), .ZN(\ML_int[9][53] ) );
  NR2D0BWP U384 ( .A1(n2), .A2(n108), .ZN(\ML_int[9][52] ) );
  NR2D0BWP U385 ( .A1(n2), .A2(n109), .ZN(\ML_int[9][51] ) );
  NR2D0BWP U386 ( .A1(n2), .A2(n110), .ZN(\ML_int[9][50] ) );
  NR2D0BWP U387 ( .A1(n2), .A2(n111), .ZN(\ML_int[9][4] ) );
  NR2D0BWP U388 ( .A1(n2), .A2(n112), .ZN(\ML_int[9][49] ) );
  NR2D0BWP U389 ( .A1(n2), .A2(n113), .ZN(\ML_int[9][48] ) );
  NR2D0BWP U390 ( .A1(n2), .A2(n114), .ZN(\ML_int[9][47] ) );
  NR2D0BWP U391 ( .A1(n2), .A2(n115), .ZN(\ML_int[9][46] ) );
  NR2D0BWP U392 ( .A1(n3), .A2(n116), .ZN(\ML_int[9][45] ) );
  NR2D0BWP U393 ( .A1(n3), .A2(n117), .ZN(\ML_int[9][44] ) );
  NR2D0BWP U394 ( .A1(n3), .A2(n118), .ZN(\ML_int[9][43] ) );
  NR2D0BWP U395 ( .A1(n3), .A2(n119), .ZN(\ML_int[9][42] ) );
  NR2D0BWP U396 ( .A1(n3), .A2(n120), .ZN(\ML_int[9][41] ) );
  NR2D0BWP U397 ( .A1(n3), .A2(n121), .ZN(\ML_int[9][40] ) );
  NR2D0BWP U398 ( .A1(n3), .A2(n122), .ZN(\ML_int[9][3] ) );
  NR2D0BWP U399 ( .A1(n3), .A2(n123), .ZN(\ML_int[9][39] ) );
  NR2D0BWP U400 ( .A1(n3), .A2(n124), .ZN(\ML_int[9][38] ) );
  NR2D0BWP U401 ( .A1(n3), .A2(n125), .ZN(\ML_int[9][37] ) );
  NR2D0BWP U402 ( .A1(n3), .A2(n126), .ZN(\ML_int[9][36] ) );
  NR2D0BWP U403 ( .A1(n3), .A2(n127), .ZN(\ML_int[9][35] ) );
  NR2D0BWP U404 ( .A1(n4), .A2(n128), .ZN(\ML_int[9][34] ) );
  NR2D0BWP U405 ( .A1(n4), .A2(n129), .ZN(\ML_int[9][33] ) );
  NR2D0BWP U406 ( .A1(n4), .A2(n130), .ZN(\ML_int[9][32] ) );
  NR2D0BWP U407 ( .A1(n4), .A2(n131), .ZN(\ML_int[9][31] ) );
  NR2D0BWP U408 ( .A1(n4), .A2(n132), .ZN(\ML_int[9][30] ) );
  NR2D0BWP U409 ( .A1(n4), .A2(n133), .ZN(\ML_int[9][2] ) );
  NR2D0BWP U410 ( .A1(n4), .A2(n134), .ZN(\ML_int[9][29] ) );
  NR2D0BWP U411 ( .A1(n4), .A2(n135), .ZN(\ML_int[9][28] ) );
  NR2D0BWP U412 ( .A1(n4), .A2(n136), .ZN(\ML_int[9][27] ) );
  NR2D0BWP U413 ( .A1(n4), .A2(n137), .ZN(\ML_int[9][26] ) );
  NR2D0BWP U414 ( .A1(n4), .A2(n138), .ZN(\ML_int[9][25] ) );
  INR2D0BWP U415 ( .A1(\ML_int[8][255] ), .B1(SH[8]), .ZN(\ML_int[9][255] ) );
  INR2D0BWP U416 ( .A1(\ML_int[8][254] ), .B1(SH[8]), .ZN(\ML_int[9][254] ) );
  INR2D0BWP U417 ( .A1(\ML_int[8][253] ), .B1(SH[8]), .ZN(\ML_int[9][253] ) );
  INR2D0BWP U418 ( .A1(\ML_int[8][252] ), .B1(SH[8]), .ZN(\ML_int[9][252] ) );
  INR2D0BWP U419 ( .A1(\ML_int[8][251] ), .B1(SH[8]), .ZN(\ML_int[9][251] ) );
  INR2D0BWP U420 ( .A1(\ML_int[8][250] ), .B1(SH[8]), .ZN(\ML_int[9][250] ) );
  NR2D0BWP U421 ( .A1(n5), .A2(n139), .ZN(\ML_int[9][24] ) );
  INR2D0BWP U422 ( .A1(\ML_int[8][249] ), .B1(SH[8]), .ZN(\ML_int[9][249] ) );
  INR2D0BWP U423 ( .A1(\ML_int[8][248] ), .B1(SH[8]), .ZN(\ML_int[9][248] ) );
  INR2D0BWP U424 ( .A1(\ML_int[8][247] ), .B1(SH[8]), .ZN(\ML_int[9][247] ) );
  INR2D0BWP U425 ( .A1(\ML_int[8][246] ), .B1(SH[8]), .ZN(\ML_int[9][246] ) );
  INR2D0BWP U426 ( .A1(\ML_int[8][245] ), .B1(SH[8]), .ZN(\ML_int[9][245] ) );
  INR2D0BWP U427 ( .A1(\ML_int[8][244] ), .B1(SH[8]), .ZN(\ML_int[9][244] ) );
  INR2D0BWP U428 ( .A1(\ML_int[8][243] ), .B1(SH[8]), .ZN(\ML_int[9][243] ) );
  INR2D0BWP U429 ( .A1(\ML_int[8][242] ), .B1(SH[8]), .ZN(\ML_int[9][242] ) );
  INR2D0BWP U430 ( .A1(\ML_int[8][241] ), .B1(SH[8]), .ZN(\ML_int[9][241] ) );
  INR2D0BWP U431 ( .A1(\ML_int[8][240] ), .B1(SH[8]), .ZN(\ML_int[9][240] ) );
  NR2D0BWP U432 ( .A1(n5), .A2(n140), .ZN(\ML_int[9][23] ) );
  INR2D0BWP U433 ( .A1(\ML_int[8][239] ), .B1(SH[8]), .ZN(\ML_int[9][239] ) );
  INR2D0BWP U434 ( .A1(\ML_int[8][238] ), .B1(SH[8]), .ZN(\ML_int[9][238] ) );
  INR2D0BWP U435 ( .A1(\ML_int[8][237] ), .B1(SH[8]), .ZN(\ML_int[9][237] ) );
  INR2D0BWP U436 ( .A1(\ML_int[8][236] ), .B1(SH[8]), .ZN(\ML_int[9][236] ) );
  INR2D0BWP U437 ( .A1(\ML_int[8][235] ), .B1(SH[8]), .ZN(\ML_int[9][235] ) );
  INR2D0BWP U438 ( .A1(\ML_int[8][234] ), .B1(SH[8]), .ZN(\ML_int[9][234] ) );
  INR2D0BWP U439 ( .A1(\ML_int[8][233] ), .B1(SH[8]), .ZN(\ML_int[9][233] ) );
  INR2D0BWP U440 ( .A1(\ML_int[8][232] ), .B1(SH[8]), .ZN(\ML_int[9][232] ) );
  INR2D0BWP U441 ( .A1(\ML_int[8][231] ), .B1(SH[8]), .ZN(\ML_int[9][231] ) );
  INR2D0BWP U442 ( .A1(\ML_int[8][230] ), .B1(SH[8]), .ZN(\ML_int[9][230] ) );
  NR2D0BWP U443 ( .A1(n5), .A2(n141), .ZN(\ML_int[9][22] ) );
  INR2D0BWP U444 ( .A1(\ML_int[8][229] ), .B1(SH[8]), .ZN(\ML_int[9][229] ) );
  INR2D0BWP U445 ( .A1(\ML_int[8][228] ), .B1(SH[8]), .ZN(\ML_int[9][228] ) );
  INR2D0BWP U446 ( .A1(\ML_int[8][227] ), .B1(SH[8]), .ZN(\ML_int[9][227] ) );
  INR2D0BWP U447 ( .A1(\ML_int[8][226] ), .B1(SH[8]), .ZN(\ML_int[9][226] ) );
  INR2D0BWP U448 ( .A1(\ML_int[8][225] ), .B1(SH[8]), .ZN(\ML_int[9][225] ) );
  INR2D0BWP U449 ( .A1(\ML_int[8][224] ), .B1(SH[8]), .ZN(\ML_int[9][224] ) );
  INR2D0BWP U450 ( .A1(\ML_int[8][223] ), .B1(SH[8]), .ZN(\ML_int[9][223] ) );
  INR2D0BWP U451 ( .A1(\ML_int[8][222] ), .B1(SH[8]), .ZN(\ML_int[9][222] ) );
  INR2D0BWP U452 ( .A1(\ML_int[8][221] ), .B1(SH[8]), .ZN(\ML_int[9][221] ) );
  INR2D0BWP U453 ( .A1(\ML_int[8][220] ), .B1(SH[8]), .ZN(\ML_int[9][220] ) );
  NR2D0BWP U454 ( .A1(n5), .A2(n142), .ZN(\ML_int[9][21] ) );
  INR2D0BWP U455 ( .A1(\ML_int[8][219] ), .B1(SH[8]), .ZN(\ML_int[9][219] ) );
  INR2D0BWP U456 ( .A1(\ML_int[8][218] ), .B1(SH[8]), .ZN(\ML_int[9][218] ) );
  INR2D0BWP U457 ( .A1(\ML_int[8][217] ), .B1(SH[8]), .ZN(\ML_int[9][217] ) );
  INR2D0BWP U458 ( .A1(\ML_int[8][216] ), .B1(SH[8]), .ZN(\ML_int[9][216] ) );
  INR2D0BWP U459 ( .A1(\ML_int[8][215] ), .B1(SH[8]), .ZN(\ML_int[9][215] ) );
  INR2D0BWP U460 ( .A1(\ML_int[8][214] ), .B1(SH[8]), .ZN(\ML_int[9][214] ) );
  INR2D0BWP U461 ( .A1(\ML_int[8][213] ), .B1(SH[8]), .ZN(\ML_int[9][213] ) );
  INR2D0BWP U462 ( .A1(\ML_int[8][212] ), .B1(SH[8]), .ZN(\ML_int[9][212] ) );
  INR2D0BWP U463 ( .A1(\ML_int[8][211] ), .B1(SH[8]), .ZN(\ML_int[9][211] ) );
  INR2D0BWP U464 ( .A1(\ML_int[8][210] ), .B1(SH[8]), .ZN(\ML_int[9][210] ) );
  NR2D0BWP U465 ( .A1(n5), .A2(n143), .ZN(\ML_int[9][20] ) );
  INR2D0BWP U466 ( .A1(\ML_int[8][209] ), .B1(SH[8]), .ZN(\ML_int[9][209] ) );
  INR2D0BWP U467 ( .A1(\ML_int[8][208] ), .B1(SH[8]), .ZN(\ML_int[9][208] ) );
  INR2D0BWP U468 ( .A1(\ML_int[8][207] ), .B1(SH[8]), .ZN(\ML_int[9][207] ) );
  INR2D0BWP U469 ( .A1(\ML_int[8][206] ), .B1(SH[8]), .ZN(\ML_int[9][206] ) );
  INR2D0BWP U470 ( .A1(\ML_int[8][205] ), .B1(SH[8]), .ZN(\ML_int[9][205] ) );
  INR2D0BWP U471 ( .A1(\ML_int[8][204] ), .B1(SH[8]), .ZN(\ML_int[9][204] ) );
  INR2D0BWP U472 ( .A1(\ML_int[8][203] ), .B1(SH[8]), .ZN(\ML_int[9][203] ) );
  INR2D0BWP U473 ( .A1(\ML_int[8][202] ), .B1(SH[8]), .ZN(\ML_int[9][202] ) );
  INR2D0BWP U474 ( .A1(\ML_int[8][201] ), .B1(SH[8]), .ZN(\ML_int[9][201] ) );
  INR2D0BWP U475 ( .A1(\ML_int[8][200] ), .B1(SH[8]), .ZN(\ML_int[9][200] ) );
  NR2D0BWP U476 ( .A1(n5), .A2(n144), .ZN(\ML_int[9][1] ) );
  NR2D0BWP U477 ( .A1(n5), .A2(n145), .ZN(\ML_int[9][19] ) );
  INR2D0BWP U478 ( .A1(\ML_int[8][199] ), .B1(SH[8]), .ZN(\ML_int[9][199] ) );
  INR2D0BWP U479 ( .A1(\ML_int[8][198] ), .B1(SH[8]), .ZN(\ML_int[9][198] ) );
  INR2D0BWP U480 ( .A1(\ML_int[8][197] ), .B1(SH[8]), .ZN(\ML_int[9][197] ) );
  INR2D0BWP U481 ( .A1(\ML_int[8][196] ), .B1(SH[8]), .ZN(\ML_int[9][196] ) );
  INR2D0BWP U482 ( .A1(\ML_int[8][195] ), .B1(SH[8]), .ZN(\ML_int[9][195] ) );
  INR2D0BWP U483 ( .A1(\ML_int[8][194] ), .B1(SH[8]), .ZN(\ML_int[9][194] ) );
  INR2D0BWP U484 ( .A1(\ML_int[8][193] ), .B1(SH[8]), .ZN(\ML_int[9][193] ) );
  INR2D0BWP U485 ( .A1(\ML_int[8][192] ), .B1(SH[8]), .ZN(\ML_int[9][192] ) );
  INR2D0BWP U486 ( .A1(\ML_int[8][191] ), .B1(SH[8]), .ZN(\ML_int[9][191] ) );
  INR2D0BWP U487 ( .A1(\ML_int[8][190] ), .B1(SH[8]), .ZN(\ML_int[9][190] ) );
  NR2D0BWP U488 ( .A1(n5), .A2(n146), .ZN(\ML_int[9][18] ) );
  INR2D0BWP U489 ( .A1(\ML_int[8][189] ), .B1(SH[8]), .ZN(\ML_int[9][189] ) );
  INR2D0BWP U490 ( .A1(\ML_int[8][188] ), .B1(SH[8]), .ZN(\ML_int[9][188] ) );
  INR2D0BWP U491 ( .A1(\ML_int[8][187] ), .B1(SH[8]), .ZN(\ML_int[9][187] ) );
  INR2D0BWP U492 ( .A1(\ML_int[8][186] ), .B1(SH[8]), .ZN(\ML_int[9][186] ) );
  INR2D0BWP U493 ( .A1(\ML_int[8][185] ), .B1(SH[8]), .ZN(\ML_int[9][185] ) );
  INR2D0BWP U494 ( .A1(\ML_int[8][184] ), .B1(SH[8]), .ZN(\ML_int[9][184] ) );
  INR2D0BWP U495 ( .A1(\ML_int[8][183] ), .B1(SH[8]), .ZN(\ML_int[9][183] ) );
  INR2D0BWP U496 ( .A1(\ML_int[8][182] ), .B1(SH[8]), .ZN(\ML_int[9][182] ) );
  INR2D0BWP U497 ( .A1(\ML_int[8][181] ), .B1(SH[8]), .ZN(\ML_int[9][181] ) );
  INR2D0BWP U498 ( .A1(\ML_int[8][180] ), .B1(SH[8]), .ZN(\ML_int[9][180] ) );
  NR2D0BWP U499 ( .A1(n5), .A2(n147), .ZN(\ML_int[9][17] ) );
  INR2D0BWP U500 ( .A1(\ML_int[8][179] ), .B1(SH[8]), .ZN(\ML_int[9][179] ) );
  INR2D0BWP U501 ( .A1(\ML_int[8][178] ), .B1(SH[8]), .ZN(\ML_int[9][178] ) );
  INR2D0BWP U502 ( .A1(\ML_int[8][177] ), .B1(SH[8]), .ZN(\ML_int[9][177] ) );
  INR2D0BWP U503 ( .A1(\ML_int[8][176] ), .B1(SH[8]), .ZN(\ML_int[9][176] ) );
  INR2D0BWP U504 ( .A1(\ML_int[8][175] ), .B1(SH[8]), .ZN(\ML_int[9][175] ) );
  INR2D0BWP U505 ( .A1(\ML_int[8][174] ), .B1(SH[8]), .ZN(\ML_int[9][174] ) );
  INR2D0BWP U506 ( .A1(\ML_int[8][173] ), .B1(SH[8]), .ZN(\ML_int[9][173] ) );
  INR2D0BWP U507 ( .A1(\ML_int[8][172] ), .B1(SH[8]), .ZN(\ML_int[9][172] ) );
  INR2D0BWP U508 ( .A1(\ML_int[8][171] ), .B1(SH[8]), .ZN(\ML_int[9][171] ) );
  INR2D0BWP U509 ( .A1(\ML_int[8][170] ), .B1(SH[8]), .ZN(\ML_int[9][170] ) );
  NR2D0BWP U510 ( .A1(n5), .A2(n148), .ZN(\ML_int[9][16] ) );
  INR2D0BWP U511 ( .A1(\ML_int[8][169] ), .B1(SH[8]), .ZN(\ML_int[9][169] ) );
  INR2D0BWP U512 ( .A1(\ML_int[8][168] ), .B1(SH[8]), .ZN(\ML_int[9][168] ) );
  INR2D0BWP U513 ( .A1(\ML_int[8][167] ), .B1(SH[8]), .ZN(\ML_int[9][167] ) );
  INR2D0BWP U514 ( .A1(\ML_int[8][166] ), .B1(SH[8]), .ZN(\ML_int[9][166] ) );
  INR2D0BWP U515 ( .A1(\ML_int[8][165] ), .B1(SH[8]), .ZN(\ML_int[9][165] ) );
  INR2D0BWP U516 ( .A1(\ML_int[8][164] ), .B1(SH[8]), .ZN(\ML_int[9][164] ) );
  INR2D0BWP U517 ( .A1(\ML_int[8][163] ), .B1(SH[8]), .ZN(\ML_int[9][163] ) );
  INR2D0BWP U518 ( .A1(\ML_int[8][162] ), .B1(SH[8]), .ZN(\ML_int[9][162] ) );
  INR2D0BWP U519 ( .A1(\ML_int[8][161] ), .B1(SH[8]), .ZN(\ML_int[9][161] ) );
  INR2D0BWP U520 ( .A1(\ML_int[8][160] ), .B1(SH[8]), .ZN(\ML_int[9][160] ) );
  NR2D0BWP U521 ( .A1(n5), .A2(n149), .ZN(\ML_int[9][15] ) );
  INR2D0BWP U522 ( .A1(\ML_int[8][159] ), .B1(SH[8]), .ZN(\ML_int[9][159] ) );
  INR2D0BWP U523 ( .A1(\ML_int[8][158] ), .B1(SH[8]), .ZN(\ML_int[9][158] ) );
  INR2D0BWP U524 ( .A1(\ML_int[8][157] ), .B1(SH[8]), .ZN(\ML_int[9][157] ) );
  INR2D0BWP U525 ( .A1(\ML_int[8][156] ), .B1(SH[8]), .ZN(\ML_int[9][156] ) );
  INR2D0BWP U526 ( .A1(\ML_int[8][155] ), .B1(SH[8]), .ZN(\ML_int[9][155] ) );
  INR2D0BWP U527 ( .A1(\ML_int[8][154] ), .B1(SH[8]), .ZN(\ML_int[9][154] ) );
  INR2D0BWP U528 ( .A1(\ML_int[8][153] ), .B1(SH[8]), .ZN(\ML_int[9][153] ) );
  INR2D0BWP U529 ( .A1(\ML_int[8][152] ), .B1(SH[8]), .ZN(\ML_int[9][152] ) );
  INR2D0BWP U530 ( .A1(\ML_int[8][151] ), .B1(SH[8]), .ZN(\ML_int[9][151] ) );
  INR2D0BWP U531 ( .A1(\ML_int[8][150] ), .B1(SH[8]), .ZN(\ML_int[9][150] ) );
  NR2D0BWP U532 ( .A1(n5), .A2(n150), .ZN(\ML_int[9][14] ) );
  INR2D0BWP U533 ( .A1(\ML_int[8][149] ), .B1(SH[8]), .ZN(\ML_int[9][149] ) );
  INR2D0BWP U534 ( .A1(\ML_int[8][148] ), .B1(SH[8]), .ZN(\ML_int[9][148] ) );
  INR2D0BWP U535 ( .A1(\ML_int[8][147] ), .B1(SH[8]), .ZN(\ML_int[9][147] ) );
  INR2D0BWP U536 ( .A1(\ML_int[8][146] ), .B1(SH[8]), .ZN(\ML_int[9][146] ) );
  INR2D0BWP U537 ( .A1(\ML_int[8][145] ), .B1(SH[8]), .ZN(\ML_int[9][145] ) );
  INR2D0BWP U538 ( .A1(\ML_int[8][144] ), .B1(SH[8]), .ZN(\ML_int[9][144] ) );
  INR2D0BWP U539 ( .A1(\ML_int[8][143] ), .B1(SH[8]), .ZN(\ML_int[9][143] ) );
  INR2D0BWP U540 ( .A1(\ML_int[8][142] ), .B1(SH[8]), .ZN(\ML_int[9][142] ) );
  INR2D0BWP U541 ( .A1(\ML_int[8][141] ), .B1(SH[8]), .ZN(\ML_int[9][141] ) );
  INR2D0BWP U542 ( .A1(\ML_int[8][140] ), .B1(SH[8]), .ZN(\ML_int[9][140] ) );
  NR2D0BWP U543 ( .A1(n6), .A2(n151), .ZN(\ML_int[9][13] ) );
  INR2D0BWP U544 ( .A1(\ML_int[8][139] ), .B1(SH[8]), .ZN(\ML_int[9][139] ) );
  INR2D0BWP U545 ( .A1(\ML_int[8][138] ), .B1(SH[8]), .ZN(\ML_int[9][138] ) );
  INR2D0BWP U546 ( .A1(\ML_int[8][137] ), .B1(SH[8]), .ZN(\ML_int[9][137] ) );
  INR2D0BWP U547 ( .A1(\ML_int[8][136] ), .B1(SH[8]), .ZN(\ML_int[9][136] ) );
  INR2D0BWP U548 ( .A1(\ML_int[8][135] ), .B1(SH[8]), .ZN(\ML_int[9][135] ) );
  INR2D0BWP U549 ( .A1(\ML_int[8][134] ), .B1(SH[8]), .ZN(\ML_int[9][134] ) );
  INR2D0BWP U550 ( .A1(\ML_int[8][133] ), .B1(SH[8]), .ZN(\ML_int[9][133] ) );
  INR2D0BWP U551 ( .A1(\ML_int[8][132] ), .B1(SH[8]), .ZN(\ML_int[9][132] ) );
  INR2D0BWP U552 ( .A1(\ML_int[8][131] ), .B1(SH[8]), .ZN(\ML_int[9][131] ) );
  INR2D0BWP U553 ( .A1(\ML_int[8][130] ), .B1(SH[8]), .ZN(\ML_int[9][130] ) );
  NR2D0BWP U554 ( .A1(n6), .A2(n152), .ZN(\ML_int[9][12] ) );
  INR2D0BWP U555 ( .A1(\ML_int[8][129] ), .B1(SH[8]), .ZN(\ML_int[9][129] ) );
  INR2D0BWP U556 ( .A1(\ML_int[8][128] ), .B1(SH[8]), .ZN(\ML_int[9][128] ) );
  INR2D0BWP U557 ( .A1(\ML_int[7][127] ), .B1(n6), .ZN(\ML_int[9][127] ) );
  INR2D0BWP U558 ( .A1(\ML_int[7][126] ), .B1(n6), .ZN(\ML_int[9][126] ) );
  INR2D0BWP U559 ( .A1(\ML_int[7][125] ), .B1(n6), .ZN(\ML_int[9][125] ) );
  INR2D0BWP U560 ( .A1(\ML_int[7][124] ), .B1(n6), .ZN(\ML_int[9][124] ) );
  INR2D0BWP U561 ( .A1(\ML_int[7][123] ), .B1(n6), .ZN(\ML_int[9][123] ) );
  INR2D0BWP U562 ( .A1(\ML_int[7][122] ), .B1(n6), .ZN(\ML_int[9][122] ) );
  INR2D0BWP U563 ( .A1(\ML_int[7][121] ), .B1(n6), .ZN(\ML_int[9][121] ) );
  INR2D0BWP U564 ( .A1(\ML_int[7][120] ), .B1(n6), .ZN(\ML_int[9][120] ) );
  NR2D0BWP U565 ( .A1(n6), .A2(n153), .ZN(\ML_int[9][11] ) );
  INR2D0BWP U566 ( .A1(\ML_int[7][119] ), .B1(n6), .ZN(\ML_int[9][119] ) );
  INR2D0BWP U567 ( .A1(\ML_int[7][118] ), .B1(n7), .ZN(\ML_int[9][118] ) );
  INR2D0BWP U568 ( .A1(\ML_int[7][117] ), .B1(n7), .ZN(\ML_int[9][117] ) );
  INR2D0BWP U569 ( .A1(\ML_int[7][116] ), .B1(n7), .ZN(\ML_int[9][116] ) );
  INR2D0BWP U570 ( .A1(\ML_int[7][115] ), .B1(n7), .ZN(\ML_int[9][115] ) );
  INR2D0BWP U571 ( .A1(\ML_int[7][114] ), .B1(n7), .ZN(\ML_int[9][114] ) );
  INR2D0BWP U572 ( .A1(\ML_int[7][113] ), .B1(n7), .ZN(\ML_int[9][113] ) );
  INR2D0BWP U573 ( .A1(\ML_int[7][112] ), .B1(n7), .ZN(\ML_int[9][112] ) );
  INR2D0BWP U574 ( .A1(\ML_int[7][111] ), .B1(n7), .ZN(\ML_int[9][111] ) );
  INR2D0BWP U575 ( .A1(\ML_int[7][110] ), .B1(n7), .ZN(\ML_int[9][110] ) );
  NR2D0BWP U576 ( .A1(n6), .A2(n154), .ZN(\ML_int[9][10] ) );
  INR2D0BWP U577 ( .A1(\ML_int[7][109] ), .B1(n7), .ZN(\ML_int[9][109] ) );
  INR2D0BWP U578 ( .A1(\ML_int[7][108] ), .B1(n7), .ZN(\ML_int[9][108] ) );
  INR2D0BWP U579 ( .A1(\ML_int[7][107] ), .B1(n7), .ZN(\ML_int[9][107] ) );
  INR2D0BWP U580 ( .A1(\ML_int[7][106] ), .B1(n7), .ZN(\ML_int[9][106] ) );
  INR2D0BWP U581 ( .A1(\ML_int[7][105] ), .B1(n8), .ZN(\ML_int[9][105] ) );
  INR2D0BWP U582 ( .A1(\ML_int[7][104] ), .B1(n8), .ZN(\ML_int[9][104] ) );
  INR2D0BWP U583 ( .A1(\ML_int[7][103] ), .B1(n8), .ZN(\ML_int[9][103] ) );
  INR2D0BWP U584 ( .A1(\ML_int[7][102] ), .B1(n9), .ZN(\ML_int[9][102] ) );
  INR2D0BWP U585 ( .A1(\ML_int[7][101] ), .B1(n10), .ZN(\ML_int[9][101] ) );
  INR2D0BWP U586 ( .A1(\ML_int[7][100] ), .B1(n11), .ZN(\ML_int[9][100] ) );
  NR2D0BWP U587 ( .A1(n4), .A2(n155), .ZN(\ML_int[9][0] ) );
  IND2D0BWP U588 ( .A1(SH[8]), .B1(n19), .ZN(n91) );
  CKND2D0BWP U589 ( .A1(\ML_int[6][9] ), .A2(n90), .ZN(n92) );
  CKND2D0BWP U590 ( .A1(\ML_int[6][8] ), .A2(n90), .ZN(n93) );
  CKND2D0BWP U591 ( .A1(\ML_int[6][7] ), .A2(n90), .ZN(n94) );
  CKND2D0BWP U592 ( .A1(\ML_int[6][6] ), .A2(n90), .ZN(n95) );
  CKND2D0BWP U593 ( .A1(\ML_int[6][63] ), .A2(n90), .ZN(n96) );
  CKND2D0BWP U594 ( .A1(\ML_int[6][62] ), .A2(n90), .ZN(n97) );
  CKND2D0BWP U595 ( .A1(\ML_int[6][61] ), .A2(n90), .ZN(n98) );
  CKND2D0BWP U596 ( .A1(\ML_int[6][60] ), .A2(n90), .ZN(n99) );
  CKND2D0BWP U597 ( .A1(\ML_int[6][5] ), .A2(n90), .ZN(n100) );
  CKND2D0BWP U598 ( .A1(\ML_int[6][59] ), .A2(n90), .ZN(n101) );
  CKND2D0BWP U599 ( .A1(\ML_int[6][58] ), .A2(n90), .ZN(n102) );
  CKND2D0BWP U600 ( .A1(\ML_int[6][57] ), .A2(n90), .ZN(n103) );
  CKND2D0BWP U601 ( .A1(\ML_int[6][56] ), .A2(n90), .ZN(n104) );
  CKND2D0BWP U602 ( .A1(\ML_int[6][55] ), .A2(n90), .ZN(n105) );
  CKND2D0BWP U603 ( .A1(\ML_int[6][54] ), .A2(n90), .ZN(n106) );
  CKND2D0BWP U604 ( .A1(\ML_int[6][53] ), .A2(n90), .ZN(n107) );
  CKND2D0BWP U605 ( .A1(\ML_int[6][52] ), .A2(n90), .ZN(n108) );
  CKND2D0BWP U606 ( .A1(\ML_int[6][51] ), .A2(n90), .ZN(n109) );
  CKND2D0BWP U607 ( .A1(\ML_int[6][50] ), .A2(n90), .ZN(n110) );
  CKND2D0BWP U608 ( .A1(\ML_int[6][4] ), .A2(n90), .ZN(n111) );
  CKND2D0BWP U609 ( .A1(\ML_int[6][49] ), .A2(n90), .ZN(n112) );
  CKND2D0BWP U610 ( .A1(\ML_int[6][48] ), .A2(n90), .ZN(n113) );
  CKND2D0BWP U611 ( .A1(\ML_int[6][47] ), .A2(n90), .ZN(n114) );
  CKND2D0BWP U612 ( .A1(\ML_int[6][46] ), .A2(n90), .ZN(n115) );
  CKND2D0BWP U613 ( .A1(\ML_int[6][45] ), .A2(n90), .ZN(n116) );
  CKND2D0BWP U614 ( .A1(\ML_int[6][44] ), .A2(n90), .ZN(n117) );
  CKND2D0BWP U615 ( .A1(\ML_int[6][43] ), .A2(n90), .ZN(n118) );
  CKND2D0BWP U616 ( .A1(\ML_int[6][42] ), .A2(n90), .ZN(n119) );
  CKND2D0BWP U617 ( .A1(\ML_int[6][41] ), .A2(n90), .ZN(n120) );
  CKND2D0BWP U618 ( .A1(\ML_int[6][40] ), .A2(n90), .ZN(n121) );
  CKND2D0BWP U619 ( .A1(\ML_int[6][3] ), .A2(n90), .ZN(n122) );
  CKND2D0BWP U620 ( .A1(\ML_int[6][39] ), .A2(n90), .ZN(n123) );
  CKND2D0BWP U621 ( .A1(\ML_int[6][38] ), .A2(n90), .ZN(n124) );
  CKND2D0BWP U622 ( .A1(\ML_int[6][37] ), .A2(n90), .ZN(n125) );
  CKND2D0BWP U623 ( .A1(\ML_int[6][36] ), .A2(n90), .ZN(n126) );
  CKND2D0BWP U624 ( .A1(\ML_int[6][35] ), .A2(n90), .ZN(n127) );
  CKND2D0BWP U625 ( .A1(\ML_int[6][34] ), .A2(n90), .ZN(n128) );
  CKND2D0BWP U626 ( .A1(\ML_int[6][33] ), .A2(n90), .ZN(n129) );
  CKND2D0BWP U627 ( .A1(\ML_int[6][32] ), .A2(n90), .ZN(n130) );
  CKND2D0BWP U628 ( .A1(\ML_int[6][31] ), .A2(n90), .ZN(n131) );
  CKND2D0BWP U629 ( .A1(\ML_int[6][30] ), .A2(n90), .ZN(n132) );
  CKND2D0BWP U630 ( .A1(\ML_int[6][2] ), .A2(n90), .ZN(n133) );
  CKND2D0BWP U631 ( .A1(\ML_int[6][29] ), .A2(n90), .ZN(n134) );
  CKND2D0BWP U632 ( .A1(\ML_int[6][28] ), .A2(n90), .ZN(n135) );
  CKND2D0BWP U633 ( .A1(\ML_int[6][27] ), .A2(n90), .ZN(n136) );
  CKND2D0BWP U634 ( .A1(\ML_int[6][26] ), .A2(n90), .ZN(n137) );
  CKND2D0BWP U635 ( .A1(\ML_int[6][25] ), .A2(n90), .ZN(n138) );
  CKND2D0BWP U636 ( .A1(\ML_int[6][24] ), .A2(n90), .ZN(n139) );
  CKND2D0BWP U637 ( .A1(\ML_int[6][23] ), .A2(n90), .ZN(n140) );
  CKND2D0BWP U638 ( .A1(\ML_int[6][22] ), .A2(n90), .ZN(n141) );
  CKND2D0BWP U639 ( .A1(\ML_int[6][21] ), .A2(n90), .ZN(n142) );
  CKND2D0BWP U640 ( .A1(\ML_int[6][20] ), .A2(n90), .ZN(n143) );
  CKND2D0BWP U641 ( .A1(\ML_int[6][1] ), .A2(n90), .ZN(n144) );
  CKND2D0BWP U642 ( .A1(\ML_int[6][19] ), .A2(n90), .ZN(n145) );
  CKND2D0BWP U643 ( .A1(\ML_int[6][18] ), .A2(n90), .ZN(n146) );
  CKND2D0BWP U644 ( .A1(\ML_int[6][17] ), .A2(n90), .ZN(n147) );
  CKND2D0BWP U645 ( .A1(\ML_int[6][16] ), .A2(n90), .ZN(n148) );
  CKND2D0BWP U646 ( .A1(\ML_int[6][15] ), .A2(n90), .ZN(n149) );
  CKND2D0BWP U647 ( .A1(\ML_int[6][14] ), .A2(n90), .ZN(n150) );
  CKND2D0BWP U648 ( .A1(\ML_int[6][13] ), .A2(n90), .ZN(n151) );
  CKND2D0BWP U649 ( .A1(\ML_int[6][12] ), .A2(n90), .ZN(n152) );
  CKND2D0BWP U650 ( .A1(\ML_int[6][11] ), .A2(n90), .ZN(n153) );
  CKND2D0BWP U651 ( .A1(\ML_int[6][10] ), .A2(n90), .ZN(n154) );
  CKND2D0BWP U652 ( .A1(\ML_int[6][0] ), .A2(n90), .ZN(n155) );
  INR2D0BWP U653 ( .A1(\ML_int[5][9] ), .B1(SH[5]), .ZN(\ML_int[6][9] ) );
  INR2D0BWP U654 ( .A1(\ML_int[5][8] ), .B1(SH[5]), .ZN(\ML_int[6][8] ) );
  INR2D0BWP U655 ( .A1(\ML_int[5][7] ), .B1(SH[5]), .ZN(\ML_int[6][7] ) );
  INR2D0BWP U656 ( .A1(\ML_int[5][6] ), .B1(SH[5]), .ZN(\ML_int[6][6] ) );
  INR2D0BWP U657 ( .A1(\ML_int[5][5] ), .B1(SH[5]), .ZN(\ML_int[6][5] ) );
  INR2D0BWP U658 ( .A1(\ML_int[5][4] ), .B1(SH[5]), .ZN(\ML_int[6][4] ) );
  INR2D0BWP U659 ( .A1(\ML_int[5][3] ), .B1(SH[5]), .ZN(\ML_int[6][3] ) );
  INR2D0BWP U660 ( .A1(\ML_int[5][31] ), .B1(SH[5]), .ZN(\ML_int[6][31] ) );
  INR2D0BWP U661 ( .A1(\ML_int[5][30] ), .B1(SH[5]), .ZN(\ML_int[6][30] ) );
  INR2D0BWP U662 ( .A1(\ML_int[5][2] ), .B1(SH[5]), .ZN(\ML_int[6][2] ) );
  INR2D0BWP U663 ( .A1(\ML_int[5][29] ), .B1(SH[5]), .ZN(\ML_int[6][29] ) );
  INR2D0BWP U664 ( .A1(\ML_int[5][28] ), .B1(SH[5]), .ZN(\ML_int[6][28] ) );
  INR2D0BWP U665 ( .A1(\ML_int[5][27] ), .B1(SH[5]), .ZN(\ML_int[6][27] ) );
  INR2D0BWP U666 ( .A1(\ML_int[5][26] ), .B1(SH[5]), .ZN(\ML_int[6][26] ) );
  INR2D0BWP U667 ( .A1(\ML_int[5][25] ), .B1(SH[5]), .ZN(\ML_int[6][25] ) );
  INR2D0BWP U668 ( .A1(\ML_int[5][24] ), .B1(SH[5]), .ZN(\ML_int[6][24] ) );
  INR2D0BWP U669 ( .A1(\ML_int[5][23] ), .B1(SH[5]), .ZN(\ML_int[6][23] ) );
  INR2D0BWP U670 ( .A1(\ML_int[5][22] ), .B1(SH[5]), .ZN(\ML_int[6][22] ) );
  INR2D0BWP U671 ( .A1(\ML_int[5][21] ), .B1(SH[5]), .ZN(\ML_int[6][21] ) );
  INR2D0BWP U672 ( .A1(\ML_int[5][20] ), .B1(SH[5]), .ZN(\ML_int[6][20] ) );
  INR2D0BWP U673 ( .A1(\ML_int[5][1] ), .B1(SH[5]), .ZN(\ML_int[6][1] ) );
  INR2D0BWP U674 ( .A1(\ML_int[5][19] ), .B1(SH[5]), .ZN(\ML_int[6][19] ) );
  INR2D0BWP U675 ( .A1(\ML_int[5][18] ), .B1(SH[5]), .ZN(\ML_int[6][18] ) );
  INR2D0BWP U676 ( .A1(\ML_int[5][17] ), .B1(SH[5]), .ZN(\ML_int[6][17] ) );
  INR2D0BWP U677 ( .A1(\ML_int[5][16] ), .B1(SH[5]), .ZN(\ML_int[6][16] ) );
  INR2D0BWP U678 ( .A1(\ML_int[5][15] ), .B1(SH[5]), .ZN(\ML_int[6][15] ) );
  INR2D0BWP U679 ( .A1(\ML_int[5][14] ), .B1(SH[5]), .ZN(\ML_int[6][14] ) );
  INR2D0BWP U680 ( .A1(\ML_int[5][13] ), .B1(SH[5]), .ZN(\ML_int[6][13] ) );
  INR2D0BWP U681 ( .A1(\ML_int[5][12] ), .B1(SH[5]), .ZN(\ML_int[6][12] ) );
  INR2D0BWP U682 ( .A1(\ML_int[5][11] ), .B1(SH[5]), .ZN(\ML_int[6][11] ) );
  INR2D0BWP U683 ( .A1(\ML_int[5][10] ), .B1(SH[5]), .ZN(\ML_int[6][10] ) );
  INR2D0BWP U684 ( .A1(\ML_int[5][0] ), .B1(SH[5]), .ZN(\ML_int[6][0] ) );
  INR2D0BWP U685 ( .A1(\ML_int[4][9] ), .B1(SH[4]), .ZN(\ML_int[5][9] ) );
  INR2D0BWP U686 ( .A1(\ML_int[4][8] ), .B1(SH[4]), .ZN(\ML_int[5][8] ) );
  INR2D0BWP U687 ( .A1(\ML_int[4][7] ), .B1(SH[4]), .ZN(\ML_int[5][7] ) );
  INR2D0BWP U688 ( .A1(\ML_int[4][6] ), .B1(SH[4]), .ZN(\ML_int[5][6] ) );
  INR2D0BWP U689 ( .A1(\ML_int[4][5] ), .B1(SH[4]), .ZN(\ML_int[5][5] ) );
  INR2D0BWP U690 ( .A1(\ML_int[4][4] ), .B1(SH[4]), .ZN(\ML_int[5][4] ) );
  INR2D0BWP U691 ( .A1(\ML_int[4][3] ), .B1(SH[4]), .ZN(\ML_int[5][3] ) );
  INR2D0BWP U692 ( .A1(\ML_int[4][2] ), .B1(SH[4]), .ZN(\ML_int[5][2] ) );
  INR2D0BWP U693 ( .A1(\ML_int[4][1] ), .B1(SH[4]), .ZN(\ML_int[5][1] ) );
  INR2D0BWP U694 ( .A1(\MR_int[4][0] ), .B1(SH[4]), .ZN(\ML_int[5][15] ) );
  INR2D0BWP U695 ( .A1(\ML_int[4][14] ), .B1(SH[4]), .ZN(\ML_int[5][14] ) );
  INR2D0BWP U696 ( .A1(\ML_int[4][13] ), .B1(SH[4]), .ZN(\ML_int[5][13] ) );
  INR2D0BWP U697 ( .A1(\ML_int[4][12] ), .B1(SH[4]), .ZN(\ML_int[5][12] ) );
  INR2D0BWP U698 ( .A1(\ML_int[4][11] ), .B1(SH[4]), .ZN(\ML_int[5][11] ) );
  INR2D0BWP U699 ( .A1(\ML_int[4][10] ), .B1(SH[4]), .ZN(\ML_int[5][10] ) );
  INR2D0BWP U700 ( .A1(\ML_int[4][0] ), .B1(SH[4]), .ZN(\ML_int[5][0] ) );
endmodule


module CVP14_DW01_decode_1 ( A, B );
  input [4:0] A;
  output [31:0] B;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;

  INVD1BWP U2 ( .I(A[2]), .ZN(n3) );
  INVD1BWP U3 ( .I(A[0]), .ZN(n2) );
  INVD1BWP U4 ( .I(A[3]), .ZN(n1) );
  NR2D0BWP U5 ( .A1(n4), .A2(n5), .ZN(B[9]) );
  NR2D0BWP U6 ( .A1(n4), .A2(n6), .ZN(B[8]) );
  NR2D0BWP U7 ( .A1(n7), .A2(n8), .ZN(B[7]) );
  NR2D0BWP U8 ( .A1(n7), .A2(n9), .ZN(B[6]) );
  NR2D0BWP U9 ( .A1(n8), .A2(n10), .ZN(B[5]) );
  NR2D0BWP U10 ( .A1(n9), .A2(n10), .ZN(B[4]) );
  NR2D0BWP U11 ( .A1(n8), .A2(n11), .ZN(B[3]) );
  NR2D0BWP U12 ( .A1(n9), .A2(n11), .ZN(B[2]) );
  NR2D0BWP U13 ( .A1(n4), .A2(n8), .ZN(B[1]) );
  CKND2D0BWP U14 ( .A1(A[0]), .A2(n1), .ZN(n8) );
  NR2D0BWP U15 ( .A1(n6), .A2(n7), .ZN(B[14]) );
  CKND2D0BWP U16 ( .A1(A[1]), .A2(n12), .ZN(n7) );
  NR2D0BWP U17 ( .A1(n5), .A2(n10), .ZN(B[13]) );
  NR2D0BWP U18 ( .A1(n6), .A2(n10), .ZN(B[12]) );
  IND2D0BWP U19 ( .A1(A[1]), .B1(n12), .ZN(n10) );
  NR2D0BWP U20 ( .A1(n5), .A2(n11), .ZN(B[11]) );
  CKND2D0BWP U21 ( .A1(A[3]), .A2(A[0]), .ZN(n5) );
  NR2D0BWP U22 ( .A1(n6), .A2(n11), .ZN(B[10]) );
  IND3D0BWP U23 ( .A1(A[4]), .B1(n3), .B2(A[1]), .ZN(n11) );
  CKND2D0BWP U24 ( .A1(A[3]), .A2(n2), .ZN(n6) );
  NR2D0BWP U25 ( .A1(n4), .A2(n9), .ZN(B[0]) );
  CKND2D0BWP U26 ( .A1(n2), .A2(n1), .ZN(n9) );
  OR3D0BWP U27 ( .A1(n12), .A2(A[1]), .A3(A[4]), .Z(n4) );
  NR2D0BWP U28 ( .A1(n3), .A2(A[4]), .ZN(n12) );
endmodule


module CVP14_DW01_ash_2 ( A, DATA_TC, SH, SH_TC, B );
  input [255:0] A;
  input [31:0] SH;
  output [255:0] B;
  input DATA_TC, SH_TC;
  wire   \temp_int_SH[7] , \temp_int_SH[6] , \temp_int_SH[5] ,
         \temp_int_SH[4] , \ML_int[4][0] , \ML_int[5][31] , \ML_int[5][30] ,
         \ML_int[5][29] , \ML_int[5][28] , \ML_int[5][27] , \ML_int[5][26] ,
         \ML_int[5][25] , \ML_int[5][24] , \ML_int[5][23] , \ML_int[5][22] ,
         \ML_int[5][21] , \ML_int[5][20] , \ML_int[5][19] , \ML_int[5][18] ,
         \ML_int[5][17] , \ML_int[5][16] , \ML_int[5][15] , \ML_int[5][14] ,
         \ML_int[5][13] , \ML_int[5][12] , \ML_int[5][11] , \ML_int[5][10] ,
         \ML_int[5][9] , \ML_int[5][8] , \ML_int[5][7] , \ML_int[5][6] ,
         \ML_int[5][5] , \ML_int[5][4] , \ML_int[5][3] , \ML_int[5][2] ,
         \ML_int[5][1] , \ML_int[5][0] , \ML_int[6][63] , \ML_int[6][62] ,
         \ML_int[6][61] , \ML_int[6][60] , \ML_int[6][59] , \ML_int[6][58] ,
         \ML_int[6][57] , \ML_int[6][56] , \ML_int[6][55] , \ML_int[6][54] ,
         \ML_int[6][53] , \ML_int[6][52] , \ML_int[6][51] , \ML_int[6][50] ,
         \ML_int[6][49] , \ML_int[6][48] , \ML_int[6][47] , \ML_int[6][46] ,
         \ML_int[6][45] , \ML_int[6][44] , \ML_int[6][43] , \ML_int[6][42] ,
         \ML_int[6][41] , \ML_int[6][40] , \ML_int[6][39] , \ML_int[6][38] ,
         \ML_int[6][37] , \ML_int[6][36] , \ML_int[6][35] , \ML_int[6][34] ,
         \ML_int[6][33] , \ML_int[6][32] , \ML_int[6][31] , \ML_int[6][30] ,
         \ML_int[6][29] , \ML_int[6][28] , \ML_int[6][27] , \ML_int[6][26] ,
         \ML_int[6][25] , \ML_int[6][24] , \ML_int[6][23] , \ML_int[6][22] ,
         \ML_int[6][21] , \ML_int[6][20] , \ML_int[6][19] , \ML_int[6][18] ,
         \ML_int[6][17] , \ML_int[6][16] , \ML_int[6][15] , \ML_int[6][14] ,
         \ML_int[6][13] , \ML_int[6][12] , \ML_int[6][11] , \ML_int[6][10] ,
         \ML_int[6][9] , \ML_int[6][8] , \ML_int[6][7] , \ML_int[6][6] ,
         \ML_int[6][5] , \ML_int[6][4] , \ML_int[6][3] , \ML_int[6][2] ,
         \ML_int[6][1] , \ML_int[6][0] , \ML_int[7][127] , \ML_int[7][126] ,
         \ML_int[7][125] , \ML_int[7][124] , \ML_int[7][123] ,
         \ML_int[7][122] , \ML_int[7][121] , \ML_int[7][120] ,
         \ML_int[7][119] , \ML_int[7][118] , \ML_int[7][117] ,
         \ML_int[7][116] , \ML_int[7][115] , \ML_int[7][114] ,
         \ML_int[7][113] , \ML_int[7][112] , \ML_int[7][111] ,
         \ML_int[7][110] , \ML_int[7][109] , \ML_int[7][108] ,
         \ML_int[7][107] , \ML_int[7][106] , \ML_int[7][105] ,
         \ML_int[7][104] , \ML_int[7][103] , \ML_int[7][102] ,
         \ML_int[7][101] , \ML_int[7][100] , \ML_int[7][99] , \ML_int[7][98] ,
         \ML_int[7][97] , \ML_int[7][96] , \ML_int[7][95] , \ML_int[7][94] ,
         \ML_int[7][93] , \ML_int[7][92] , \ML_int[7][91] , \ML_int[7][90] ,
         \ML_int[7][89] , \ML_int[7][88] , \ML_int[7][87] , \ML_int[7][86] ,
         \ML_int[7][85] , \ML_int[7][84] , \ML_int[7][83] , \ML_int[7][82] ,
         \ML_int[7][81] , \ML_int[7][80] , \ML_int[7][79] , \ML_int[7][78] ,
         \ML_int[7][77] , \ML_int[7][76] , \ML_int[7][75] , \ML_int[7][74] ,
         \ML_int[7][73] , \ML_int[7][72] , \ML_int[7][71] , \ML_int[7][70] ,
         \ML_int[7][69] , \ML_int[7][68] , \ML_int[7][67] , \ML_int[7][66] ,
         \ML_int[7][65] , \ML_int[7][64] , \ML_int[8][255] , \ML_int[8][254] ,
         \ML_int[8][253] , \ML_int[8][252] , \ML_int[8][251] ,
         \ML_int[8][250] , \ML_int[8][249] , \ML_int[8][248] ,
         \ML_int[8][247] , \ML_int[8][246] , \ML_int[8][245] ,
         \ML_int[8][244] , \ML_int[8][243] , \ML_int[8][242] ,
         \ML_int[8][241] , \ML_int[8][240] , \ML_int[8][239] ,
         \ML_int[8][238] , \ML_int[8][237] , \ML_int[8][236] ,
         \ML_int[8][235] , \ML_int[8][234] , \ML_int[8][233] ,
         \ML_int[8][232] , \ML_int[8][231] , \ML_int[8][230] ,
         \ML_int[8][229] , \ML_int[8][228] , \ML_int[8][227] ,
         \ML_int[8][226] , \ML_int[8][225] , \ML_int[8][224] ,
         \ML_int[8][223] , \ML_int[8][222] , \ML_int[8][221] ,
         \ML_int[8][220] , \ML_int[8][219] , \ML_int[8][218] ,
         \ML_int[8][217] , \ML_int[8][216] , \ML_int[8][215] ,
         \ML_int[8][214] , \ML_int[8][213] , \ML_int[8][212] ,
         \ML_int[8][211] , \ML_int[8][210] , \ML_int[8][209] ,
         \ML_int[8][208] , \ML_int[8][207] , \ML_int[8][206] ,
         \ML_int[8][205] , \ML_int[8][204] , \ML_int[8][203] ,
         \ML_int[8][202] , \ML_int[8][201] , \ML_int[8][200] ,
         \ML_int[8][199] , \ML_int[8][198] , \ML_int[8][197] ,
         \ML_int[8][196] , \ML_int[8][195] , \ML_int[8][194] ,
         \ML_int[8][193] , \ML_int[8][192] , \ML_int[8][191] ,
         \ML_int[8][190] , \ML_int[8][189] , \ML_int[8][188] ,
         \ML_int[8][187] , \ML_int[8][186] , \ML_int[8][185] ,
         \ML_int[8][184] , \ML_int[8][183] , \ML_int[8][182] ,
         \ML_int[8][181] , \ML_int[8][180] , \ML_int[8][179] ,
         \ML_int[8][178] , \ML_int[8][177] , \ML_int[8][176] ,
         \ML_int[8][175] , \ML_int[8][174] , \ML_int[8][173] ,
         \ML_int[8][172] , \ML_int[8][171] , \ML_int[8][170] ,
         \ML_int[8][169] , \ML_int[8][168] , \ML_int[8][167] ,
         \ML_int[8][166] , \ML_int[8][165] , \ML_int[8][164] ,
         \ML_int[8][163] , \ML_int[8][162] , \ML_int[8][161] ,
         \ML_int[8][160] , \ML_int[8][159] , \ML_int[8][158] ,
         \ML_int[8][157] , \ML_int[8][156] , \ML_int[8][155] ,
         \ML_int[8][154] , \ML_int[8][153] , \ML_int[8][152] ,
         \ML_int[8][151] , \ML_int[8][150] , \ML_int[8][149] ,
         \ML_int[8][148] , \ML_int[8][147] , \ML_int[8][146] ,
         \ML_int[8][145] , \ML_int[8][144] , \ML_int[8][143] ,
         \ML_int[8][142] , \ML_int[8][141] , \ML_int[8][140] ,
         \ML_int[8][139] , \ML_int[8][138] , \ML_int[8][137] ,
         \ML_int[8][136] , \ML_int[8][135] , \ML_int[8][134] ,
         \ML_int[8][133] , \ML_int[8][132] , \ML_int[8][131] ,
         \ML_int[8][130] , \ML_int[8][129] , \ML_int[8][128] ,
         \ML_int[10][255] , \ML_int[10][254] , \ML_int[10][253] ,
         \ML_int[10][252] , \ML_int[10][251] , \ML_int[10][250] ,
         \ML_int[10][249] , \ML_int[10][248] , \ML_int[10][247] ,
         \ML_int[10][246] , \ML_int[10][245] , \ML_int[10][244] ,
         \ML_int[10][243] , \ML_int[10][242] , \ML_int[10][241] ,
         \ML_int[10][240] , \ML_int[10][239] , \ML_int[10][238] ,
         \ML_int[10][237] , \ML_int[10][236] , \ML_int[10][235] ,
         \ML_int[10][234] , \ML_int[10][233] , \ML_int[10][232] ,
         \ML_int[10][231] , \ML_int[10][230] , \ML_int[10][229] ,
         \ML_int[10][228] , \ML_int[10][227] , \ML_int[10][226] ,
         \ML_int[10][225] , \ML_int[10][224] , \ML_int[10][223] ,
         \ML_int[10][222] , \ML_int[10][221] , \ML_int[10][220] ,
         \ML_int[10][219] , \ML_int[10][218] , \ML_int[10][217] ,
         \ML_int[10][216] , \ML_int[10][215] , \ML_int[10][214] ,
         \ML_int[10][213] , \ML_int[10][212] , \ML_int[10][211] ,
         \ML_int[10][210] , \ML_int[10][209] , \ML_int[10][208] ,
         \ML_int[10][207] , \ML_int[10][206] , \ML_int[10][205] ,
         \ML_int[10][204] , \ML_int[10][203] , \ML_int[10][202] ,
         \ML_int[10][201] , \ML_int[10][200] , \ML_int[10][199] ,
         \ML_int[10][198] , \ML_int[10][197] , \ML_int[10][196] ,
         \ML_int[10][195] , \ML_int[10][194] , \ML_int[10][193] ,
         \ML_int[10][192] , \ML_int[10][191] , \ML_int[10][190] ,
         \ML_int[10][189] , \ML_int[10][188] , \ML_int[10][187] ,
         \ML_int[10][186] , \ML_int[10][185] , \ML_int[10][184] ,
         \ML_int[10][183] , \ML_int[10][182] , \ML_int[10][181] ,
         \ML_int[10][180] , \ML_int[10][179] , \ML_int[10][178] ,
         \ML_int[10][177] , \ML_int[10][176] , \ML_int[10][175] ,
         \ML_int[10][174] , \ML_int[10][173] , \ML_int[10][172] ,
         \ML_int[10][171] , \ML_int[10][170] , \ML_int[10][169] ,
         \ML_int[10][168] , \ML_int[10][167] , \ML_int[10][166] ,
         \ML_int[10][165] , \ML_int[10][164] , \ML_int[10][163] ,
         \ML_int[10][162] , \ML_int[10][161] , \ML_int[10][160] ,
         \ML_int[10][159] , \ML_int[10][158] , \ML_int[10][157] ,
         \ML_int[10][156] , \ML_int[10][155] , \ML_int[10][154] ,
         \ML_int[10][153] , \ML_int[10][152] , \ML_int[10][151] ,
         \ML_int[10][150] , \ML_int[10][149] , \ML_int[10][148] ,
         \ML_int[10][147] , \ML_int[10][146] , \ML_int[10][145] ,
         \ML_int[10][144] , \ML_int[10][143] , \ML_int[10][142] ,
         \ML_int[10][141] , \ML_int[10][140] , \ML_int[10][139] ,
         \ML_int[10][138] , \ML_int[10][137] , \ML_int[10][136] ,
         \ML_int[10][135] , \ML_int[10][134] , \ML_int[10][133] ,
         \ML_int[10][132] , \ML_int[10][131] , \ML_int[10][130] ,
         \ML_int[10][129] , \ML_int[10][128] , \ML_int[10][127] ,
         \ML_int[10][126] , \ML_int[10][125] , \ML_int[10][124] ,
         \ML_int[10][123] , \ML_int[10][122] , \ML_int[10][121] ,
         \ML_int[10][120] , \ML_int[10][119] , \ML_int[10][118] ,
         \ML_int[10][117] , \ML_int[10][116] , \ML_int[10][115] ,
         \ML_int[10][114] , \ML_int[10][113] , \ML_int[10][112] ,
         \ML_int[10][111] , \ML_int[10][110] , \ML_int[10][109] ,
         \ML_int[10][108] , \ML_int[10][107] , \ML_int[10][106] ,
         \ML_int[10][105] , \ML_int[10][104] , \ML_int[10][103] ,
         \ML_int[10][102] , \ML_int[10][101] , \ML_int[10][100] ,
         \ML_int[10][99] , \ML_int[10][98] , \ML_int[10][97] ,
         \ML_int[10][96] , \ML_int[10][95] , \ML_int[10][94] ,
         \ML_int[10][93] , \ML_int[10][92] , \ML_int[10][91] ,
         \ML_int[10][90] , \ML_int[10][89] , \ML_int[10][88] ,
         \ML_int[10][87] , \ML_int[10][86] , \ML_int[10][85] ,
         \ML_int[10][84] , \ML_int[10][83] , \ML_int[10][82] ,
         \ML_int[10][81] , \ML_int[10][80] , \ML_int[10][79] ,
         \ML_int[10][78] , \ML_int[10][77] , \ML_int[10][76] ,
         \ML_int[10][75] , \ML_int[10][74] , \ML_int[10][73] ,
         \ML_int[10][72] , \ML_int[10][71] , \ML_int[10][70] ,
         \ML_int[10][69] , \ML_int[10][68] , \ML_int[10][67] ,
         \ML_int[10][66] , \ML_int[10][65] , \ML_int[10][64] ,
         \ML_int[10][63] , \ML_int[10][62] , \ML_int[10][61] ,
         \ML_int[10][60] , \ML_int[10][59] , \ML_int[10][58] ,
         \ML_int[10][57] , \ML_int[10][56] , \ML_int[10][55] ,
         \ML_int[10][54] , \ML_int[10][53] , \ML_int[10][52] ,
         \ML_int[10][51] , \ML_int[10][50] , \ML_int[10][49] ,
         \ML_int[10][48] , \ML_int[10][47] , \ML_int[10][46] ,
         \ML_int[10][45] , \ML_int[10][44] , \ML_int[10][43] ,
         \ML_int[10][42] , \ML_int[10][41] , \ML_int[10][40] ,
         \ML_int[10][39] , \ML_int[10][38] , \ML_int[10][37] ,
         \ML_int[10][36] , \ML_int[10][35] , \ML_int[10][34] ,
         \ML_int[10][33] , \ML_int[10][32] , \ML_int[10][31] ,
         \ML_int[10][30] , \ML_int[10][29] , \ML_int[10][28] ,
         \ML_int[10][27] , \ML_int[10][26] , \ML_int[10][25] ,
         \ML_int[10][24] , \ML_int[10][23] , \ML_int[10][22] ,
         \ML_int[10][21] , \ML_int[10][20] , \ML_int[10][19] ,
         \ML_int[10][18] , \ML_int[10][17] , \ML_int[10][16] ,
         \ML_int[10][15] , \ML_int[10][14] , \ML_int[10][13] ,
         \ML_int[10][12] , \ML_int[10][11] , \ML_int[10][10] , \ML_int[10][9] ,
         \ML_int[10][8] , \ML_int[10][7] , \ML_int[10][6] , \ML_int[10][5] ,
         \ML_int[10][4] , \ML_int[10][3] , \ML_int[10][2] , \ML_int[10][1] ,
         \ML_int[10][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173;
  assign \temp_int_SH[7]  = SH[7];
  assign \temp_int_SH[6]  = SH[6];
  assign \temp_int_SH[5]  = SH[5];
  assign \temp_int_SH[4]  = SH[4];
  assign \ML_int[4][0]  = A[0];
  assign B[255] = \ML_int[10][255] ;
  assign B[254] = \ML_int[10][254] ;
  assign B[253] = \ML_int[10][253] ;
  assign B[252] = \ML_int[10][252] ;
  assign B[251] = \ML_int[10][251] ;
  assign B[250] = \ML_int[10][250] ;
  assign B[249] = \ML_int[10][249] ;
  assign B[248] = \ML_int[10][248] ;
  assign B[247] = \ML_int[10][247] ;
  assign B[246] = \ML_int[10][246] ;
  assign B[245] = \ML_int[10][245] ;
  assign B[244] = \ML_int[10][244] ;
  assign B[243] = \ML_int[10][243] ;
  assign B[242] = \ML_int[10][242] ;
  assign B[241] = \ML_int[10][241] ;
  assign B[240] = \ML_int[10][240] ;
  assign B[239] = \ML_int[10][239] ;
  assign B[238] = \ML_int[10][238] ;
  assign B[237] = \ML_int[10][237] ;
  assign B[236] = \ML_int[10][236] ;
  assign B[235] = \ML_int[10][235] ;
  assign B[234] = \ML_int[10][234] ;
  assign B[233] = \ML_int[10][233] ;
  assign B[232] = \ML_int[10][232] ;
  assign B[231] = \ML_int[10][231] ;
  assign B[230] = \ML_int[10][230] ;
  assign B[229] = \ML_int[10][229] ;
  assign B[228] = \ML_int[10][228] ;
  assign B[227] = \ML_int[10][227] ;
  assign B[226] = \ML_int[10][226] ;
  assign B[225] = \ML_int[10][225] ;
  assign B[224] = \ML_int[10][224] ;
  assign B[223] = \ML_int[10][223] ;
  assign B[222] = \ML_int[10][222] ;
  assign B[221] = \ML_int[10][221] ;
  assign B[220] = \ML_int[10][220] ;
  assign B[219] = \ML_int[10][219] ;
  assign B[218] = \ML_int[10][218] ;
  assign B[217] = \ML_int[10][217] ;
  assign B[216] = \ML_int[10][216] ;
  assign B[215] = \ML_int[10][215] ;
  assign B[214] = \ML_int[10][214] ;
  assign B[213] = \ML_int[10][213] ;
  assign B[212] = \ML_int[10][212] ;
  assign B[211] = \ML_int[10][211] ;
  assign B[210] = \ML_int[10][210] ;
  assign B[209] = \ML_int[10][209] ;
  assign B[208] = \ML_int[10][208] ;
  assign B[207] = \ML_int[10][207] ;
  assign B[206] = \ML_int[10][206] ;
  assign B[205] = \ML_int[10][205] ;
  assign B[204] = \ML_int[10][204] ;
  assign B[203] = \ML_int[10][203] ;
  assign B[202] = \ML_int[10][202] ;
  assign B[201] = \ML_int[10][201] ;
  assign B[200] = \ML_int[10][200] ;
  assign B[199] = \ML_int[10][199] ;
  assign B[198] = \ML_int[10][198] ;
  assign B[197] = \ML_int[10][197] ;
  assign B[196] = \ML_int[10][196] ;
  assign B[195] = \ML_int[10][195] ;
  assign B[194] = \ML_int[10][194] ;
  assign B[193] = \ML_int[10][193] ;
  assign B[192] = \ML_int[10][192] ;
  assign B[191] = \ML_int[10][191] ;
  assign B[190] = \ML_int[10][190] ;
  assign B[189] = \ML_int[10][189] ;
  assign B[188] = \ML_int[10][188] ;
  assign B[187] = \ML_int[10][187] ;
  assign B[186] = \ML_int[10][186] ;
  assign B[185] = \ML_int[10][185] ;
  assign B[184] = \ML_int[10][184] ;
  assign B[183] = \ML_int[10][183] ;
  assign B[182] = \ML_int[10][182] ;
  assign B[181] = \ML_int[10][181] ;
  assign B[180] = \ML_int[10][180] ;
  assign B[179] = \ML_int[10][179] ;
  assign B[178] = \ML_int[10][178] ;
  assign B[177] = \ML_int[10][177] ;
  assign B[176] = \ML_int[10][176] ;
  assign B[175] = \ML_int[10][175] ;
  assign B[174] = \ML_int[10][174] ;
  assign B[173] = \ML_int[10][173] ;
  assign B[172] = \ML_int[10][172] ;
  assign B[171] = \ML_int[10][171] ;
  assign B[170] = \ML_int[10][170] ;
  assign B[169] = \ML_int[10][169] ;
  assign B[168] = \ML_int[10][168] ;
  assign B[167] = \ML_int[10][167] ;
  assign B[166] = \ML_int[10][166] ;
  assign B[165] = \ML_int[10][165] ;
  assign B[164] = \ML_int[10][164] ;
  assign B[163] = \ML_int[10][163] ;
  assign B[162] = \ML_int[10][162] ;
  assign B[161] = \ML_int[10][161] ;
  assign B[160] = \ML_int[10][160] ;
  assign B[159] = \ML_int[10][159] ;
  assign B[158] = \ML_int[10][158] ;
  assign B[157] = \ML_int[10][157] ;
  assign B[156] = \ML_int[10][156] ;
  assign B[155] = \ML_int[10][155] ;
  assign B[154] = \ML_int[10][154] ;
  assign B[153] = \ML_int[10][153] ;
  assign B[152] = \ML_int[10][152] ;
  assign B[151] = \ML_int[10][151] ;
  assign B[150] = \ML_int[10][150] ;
  assign B[149] = \ML_int[10][149] ;
  assign B[148] = \ML_int[10][148] ;
  assign B[147] = \ML_int[10][147] ;
  assign B[146] = \ML_int[10][146] ;
  assign B[145] = \ML_int[10][145] ;
  assign B[144] = \ML_int[10][144] ;
  assign B[143] = \ML_int[10][143] ;
  assign B[142] = \ML_int[10][142] ;
  assign B[141] = \ML_int[10][141] ;
  assign B[140] = \ML_int[10][140] ;
  assign B[139] = \ML_int[10][139] ;
  assign B[138] = \ML_int[10][138] ;
  assign B[137] = \ML_int[10][137] ;
  assign B[136] = \ML_int[10][136] ;
  assign B[135] = \ML_int[10][135] ;
  assign B[134] = \ML_int[10][134] ;
  assign B[133] = \ML_int[10][133] ;
  assign B[132] = \ML_int[10][132] ;
  assign B[131] = \ML_int[10][131] ;
  assign B[130] = \ML_int[10][130] ;
  assign B[129] = \ML_int[10][129] ;
  assign B[128] = \ML_int[10][128] ;
  assign B[127] = \ML_int[10][127] ;
  assign B[126] = \ML_int[10][126] ;
  assign B[125] = \ML_int[10][125] ;
  assign B[124] = \ML_int[10][124] ;
  assign B[123] = \ML_int[10][123] ;
  assign B[122] = \ML_int[10][122] ;
  assign B[121] = \ML_int[10][121] ;
  assign B[120] = \ML_int[10][120] ;
  assign B[119] = \ML_int[10][119] ;
  assign B[118] = \ML_int[10][118] ;
  assign B[117] = \ML_int[10][117] ;
  assign B[116] = \ML_int[10][116] ;
  assign B[115] = \ML_int[10][115] ;
  assign B[114] = \ML_int[10][114] ;
  assign B[113] = \ML_int[10][113] ;
  assign B[112] = \ML_int[10][112] ;
  assign B[111] = \ML_int[10][111] ;
  assign B[110] = \ML_int[10][110] ;
  assign B[109] = \ML_int[10][109] ;
  assign B[108] = \ML_int[10][108] ;
  assign B[107] = \ML_int[10][107] ;
  assign B[106] = \ML_int[10][106] ;
  assign B[105] = \ML_int[10][105] ;
  assign B[104] = \ML_int[10][104] ;
  assign B[103] = \ML_int[10][103] ;
  assign B[102] = \ML_int[10][102] ;
  assign B[101] = \ML_int[10][101] ;
  assign B[100] = \ML_int[10][100] ;
  assign B[99] = \ML_int[10][99] ;
  assign B[98] = \ML_int[10][98] ;
  assign B[97] = \ML_int[10][97] ;
  assign B[96] = \ML_int[10][96] ;
  assign B[95] = \ML_int[10][95] ;
  assign B[94] = \ML_int[10][94] ;
  assign B[93] = \ML_int[10][93] ;
  assign B[92] = \ML_int[10][92] ;
  assign B[91] = \ML_int[10][91] ;
  assign B[90] = \ML_int[10][90] ;
  assign B[89] = \ML_int[10][89] ;
  assign B[88] = \ML_int[10][88] ;
  assign B[87] = \ML_int[10][87] ;
  assign B[86] = \ML_int[10][86] ;
  assign B[85] = \ML_int[10][85] ;
  assign B[84] = \ML_int[10][84] ;
  assign B[83] = \ML_int[10][83] ;
  assign B[82] = \ML_int[10][82] ;
  assign B[81] = \ML_int[10][81] ;
  assign B[80] = \ML_int[10][80] ;
  assign B[79] = \ML_int[10][79] ;
  assign B[78] = \ML_int[10][78] ;
  assign B[77] = \ML_int[10][77] ;
  assign B[76] = \ML_int[10][76] ;
  assign B[75] = \ML_int[10][75] ;
  assign B[74] = \ML_int[10][74] ;
  assign B[73] = \ML_int[10][73] ;
  assign B[72] = \ML_int[10][72] ;
  assign B[71] = \ML_int[10][71] ;
  assign B[70] = \ML_int[10][70] ;
  assign B[69] = \ML_int[10][69] ;
  assign B[68] = \ML_int[10][68] ;
  assign B[67] = \ML_int[10][67] ;
  assign B[66] = \ML_int[10][66] ;
  assign B[65] = \ML_int[10][65] ;
  assign B[64] = \ML_int[10][64] ;
  assign B[63] = \ML_int[10][63] ;
  assign B[62] = \ML_int[10][62] ;
  assign B[61] = \ML_int[10][61] ;
  assign B[60] = \ML_int[10][60] ;
  assign B[59] = \ML_int[10][59] ;
  assign B[58] = \ML_int[10][58] ;
  assign B[57] = \ML_int[10][57] ;
  assign B[56] = \ML_int[10][56] ;
  assign B[55] = \ML_int[10][55] ;
  assign B[54] = \ML_int[10][54] ;
  assign B[53] = \ML_int[10][53] ;
  assign B[52] = \ML_int[10][52] ;
  assign B[51] = \ML_int[10][51] ;
  assign B[50] = \ML_int[10][50] ;
  assign B[49] = \ML_int[10][49] ;
  assign B[48] = \ML_int[10][48] ;
  assign B[47] = \ML_int[10][47] ;
  assign B[46] = \ML_int[10][46] ;
  assign B[45] = \ML_int[10][45] ;
  assign B[44] = \ML_int[10][44] ;
  assign B[43] = \ML_int[10][43] ;
  assign B[42] = \ML_int[10][42] ;
  assign B[41] = \ML_int[10][41] ;
  assign B[40] = \ML_int[10][40] ;
  assign B[39] = \ML_int[10][39] ;
  assign B[38] = \ML_int[10][38] ;
  assign B[37] = \ML_int[10][37] ;
  assign B[36] = \ML_int[10][36] ;
  assign B[35] = \ML_int[10][35] ;
  assign B[34] = \ML_int[10][34] ;
  assign B[33] = \ML_int[10][33] ;
  assign B[32] = \ML_int[10][32] ;
  assign B[31] = \ML_int[10][31] ;
  assign B[30] = \ML_int[10][30] ;
  assign B[29] = \ML_int[10][29] ;
  assign B[28] = \ML_int[10][28] ;
  assign B[27] = \ML_int[10][27] ;
  assign B[26] = \ML_int[10][26] ;
  assign B[25] = \ML_int[10][25] ;
  assign B[24] = \ML_int[10][24] ;
  assign B[23] = \ML_int[10][23] ;
  assign B[22] = \ML_int[10][22] ;
  assign B[21] = \ML_int[10][21] ;
  assign B[20] = \ML_int[10][20] ;
  assign B[19] = \ML_int[10][19] ;
  assign B[18] = \ML_int[10][18] ;
  assign B[17] = \ML_int[10][17] ;
  assign B[16] = \ML_int[10][16] ;
  assign B[15] = \ML_int[10][15] ;
  assign B[14] = \ML_int[10][14] ;
  assign B[13] = \ML_int[10][13] ;
  assign B[12] = \ML_int[10][12] ;
  assign B[11] = \ML_int[10][11] ;
  assign B[10] = \ML_int[10][10] ;
  assign B[9] = \ML_int[10][9] ;
  assign B[8] = \ML_int[10][8] ;
  assign B[7] = \ML_int[10][7] ;
  assign B[6] = \ML_int[10][6] ;
  assign B[5] = \ML_int[10][5] ;
  assign B[4] = \ML_int[10][4] ;
  assign B[3] = \ML_int[10][3] ;
  assign B[2] = \ML_int[10][2] ;
  assign B[1] = \ML_int[10][1] ;
  assign B[0] = \ML_int[10][0] ;

  CKAN2D1BWP U3 ( .A1(\ML_int[6][54] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][118] ) );
  CKAN2D0BWP U4 ( .A1(\ML_int[6][53] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][117] ) );
  CKAN2D0BWP U5 ( .A1(\ML_int[6][52] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][116] ) );
  CKAN2D0BWP U6 ( .A1(\ML_int[6][51] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][115] ) );
  CKAN2D0BWP U7 ( .A1(\ML_int[6][50] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][114] ) );
  CKAN2D0BWP U8 ( .A1(\ML_int[6][49] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][113] ) );
  CKAN2D0BWP U9 ( .A1(\ML_int[6][48] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][112] ) );
  CKAN2D0BWP U10 ( .A1(\ML_int[6][47] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][111] ) );
  CKAN2D0BWP U11 ( .A1(\ML_int[6][46] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][110] ) );
  CKAN2D0BWP U12 ( .A1(\ML_int[6][45] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][109] ) );
  CKAN2D0BWP U13 ( .A1(\ML_int[6][44] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][108] ) );
  CKAN2D0BWP U14 ( .A1(\ML_int[6][43] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][107] ) );
  CKAN2D0BWP U15 ( .A1(\ML_int[6][42] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][106] ) );
  CKAN2D0BWP U16 ( .A1(\ML_int[6][41] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][105] ) );
  CKAN2D0BWP U17 ( .A1(\ML_int[6][40] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][104] ) );
  CKAN2D0BWP U18 ( .A1(\ML_int[6][39] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][103] ) );
  CKAN2D0BWP U19 ( .A1(\ML_int[6][38] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][102] ) );
  CKAN2D0BWP U20 ( .A1(\ML_int[6][37] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][101] ) );
  CKAN2D0BWP U21 ( .A1(\ML_int[6][36] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][100] ) );
  CKAN2D0BWP U22 ( .A1(\ML_int[6][35] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][99] ) );
  CKAN2D0BWP U23 ( .A1(\ML_int[6][34] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][98] ) );
  CKAN2D0BWP U24 ( .A1(\ML_int[6][33] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][97] ) );
  CKAN2D0BWP U25 ( .A1(\ML_int[6][32] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][96] ) );
  CKAN2D0BWP U26 ( .A1(\ML_int[6][31] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][95] ) );
  CKAN2D0BWP U27 ( .A1(\ML_int[6][30] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][94] ) );
  CKAN2D0BWP U28 ( .A1(\ML_int[6][29] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][93] ) );
  CKAN2D0BWP U29 ( .A1(\ML_int[6][28] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][92] ) );
  CKAN2D0BWP U30 ( .A1(\ML_int[6][27] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][91] ) );
  CKAN2D0BWP U31 ( .A1(\ML_int[6][26] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][90] ) );
  CKAN2D0BWP U32 ( .A1(\ML_int[6][25] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][89] ) );
  CKAN2D0BWP U33 ( .A1(\ML_int[6][24] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][88] ) );
  CKAN2D0BWP U34 ( .A1(\ML_int[6][23] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][87] ) );
  CKAN2D0BWP U35 ( .A1(\ML_int[6][22] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][86] ) );
  CKAN2D0BWP U36 ( .A1(\ML_int[6][21] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][85] ) );
  CKAN2D0BWP U37 ( .A1(\ML_int[6][20] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][84] ) );
  CKAN2D0BWP U38 ( .A1(\ML_int[6][19] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][83] ) );
  CKAN2D0BWP U39 ( .A1(\ML_int[6][18] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][82] ) );
  CKAN2D0BWP U40 ( .A1(\ML_int[6][17] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][81] ) );
  CKAN2D0BWP U41 ( .A1(\ML_int[6][16] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][80] ) );
  CKAN2D0BWP U42 ( .A1(\ML_int[6][15] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][79] ) );
  CKAN2D0BWP U43 ( .A1(\ML_int[6][14] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][78] ) );
  CKAN2D0BWP U44 ( .A1(\ML_int[6][13] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][77] ) );
  CKAN2D0BWP U45 ( .A1(\ML_int[6][12] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][76] ) );
  CKAN2D0BWP U46 ( .A1(\ML_int[6][11] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][75] ) );
  CKAN2D0BWP U47 ( .A1(\ML_int[6][10] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][74] ) );
  CKAN2D0BWP U48 ( .A1(\ML_int[6][9] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][73] ) );
  CKAN2D0BWP U49 ( .A1(\ML_int[6][8] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][72] ) );
  CKAN2D0BWP U50 ( .A1(\ML_int[6][7] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][71] ) );
  CKAN2D0BWP U51 ( .A1(\ML_int[6][6] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][70] ) );
  CKAN2D0BWP U52 ( .A1(\ML_int[6][5] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][69] ) );
  CKAN2D0BWP U53 ( .A1(\ML_int[6][4] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][68] ) );
  CKAN2D0BWP U54 ( .A1(\ML_int[6][3] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][67] ) );
  CKAN2D0BWP U55 ( .A1(\ML_int[6][2] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][66] ) );
  CKAN2D0BWP U56 ( .A1(\ML_int[6][1] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][65] ) );
  CKAN2D0BWP U57 ( .A1(\ML_int[6][0] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][64] ) );
  CKAN2D0BWP U58 ( .A1(\ML_int[5][31] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][63] ) );
  CKAN2D0BWP U59 ( .A1(\ML_int[5][30] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][62] ) );
  CKAN2D0BWP U60 ( .A1(\ML_int[5][29] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][61] ) );
  CKAN2D0BWP U61 ( .A1(\ML_int[5][28] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][60] ) );
  CKAN2D0BWP U62 ( .A1(\ML_int[5][27] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][59] ) );
  CKAN2D0BWP U63 ( .A1(\ML_int[5][26] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][58] ) );
  CKAN2D0BWP U64 ( .A1(\ML_int[5][25] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][57] ) );
  CKAN2D0BWP U65 ( .A1(\ML_int[5][24] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][56] ) );
  CKAN2D0BWP U66 ( .A1(\ML_int[5][23] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][55] ) );
  CKAN2D0BWP U67 ( .A1(\ML_int[5][22] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][54] ) );
  CKAN2D0BWP U68 ( .A1(\ML_int[5][21] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][53] ) );
  CKAN2D0BWP U69 ( .A1(\ML_int[5][20] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][52] ) );
  CKAN2D0BWP U70 ( .A1(\ML_int[5][19] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][51] ) );
  CKAN2D0BWP U71 ( .A1(\ML_int[5][18] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][50] ) );
  CKAN2D0BWP U72 ( .A1(\ML_int[5][17] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][49] ) );
  CKAN2D0BWP U73 ( .A1(\ML_int[5][16] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][48] ) );
  CKAN2D0BWP U74 ( .A1(\ML_int[5][15] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][47] ) );
  CKAN2D0BWP U75 ( .A1(\ML_int[5][14] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][46] ) );
  CKAN2D0BWP U76 ( .A1(\ML_int[5][13] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][45] ) );
  CKAN2D0BWP U77 ( .A1(\ML_int[5][12] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][44] ) );
  CKAN2D0BWP U78 ( .A1(\ML_int[5][11] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][43] ) );
  CKAN2D0BWP U79 ( .A1(\ML_int[5][10] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][42] ) );
  CKAN2D0BWP U80 ( .A1(\ML_int[5][9] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][41] ) );
  CKAN2D0BWP U81 ( .A1(\ML_int[5][8] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][40] ) );
  CKAN2D0BWP U82 ( .A1(\ML_int[5][7] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][39] ) );
  CKAN2D0BWP U83 ( .A1(\ML_int[5][6] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][38] ) );
  CKAN2D0BWP U84 ( .A1(\ML_int[5][5] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][37] ) );
  CKAN2D0BWP U85 ( .A1(\ML_int[5][4] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][36] ) );
  CKAN2D0BWP U86 ( .A1(\ML_int[5][3] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][35] ) );
  CKAN2D0BWP U87 ( .A1(\ML_int[5][2] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][34] ) );
  CKAN2D0BWP U88 ( .A1(\ML_int[5][1] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][33] ) );
  CKAN2D0BWP U89 ( .A1(\ML_int[5][0] ), .A2(\temp_int_SH[5] ), .Z(
        \ML_int[6][32] ) );
  CKBD1BWP U90 ( .I(n13), .Z(n6) );
  CKBD1BWP U91 ( .I(n13), .Z(n7) );
  CKBD1BWP U92 ( .I(n12), .Z(n10) );
  CKBD1BWP U93 ( .I(n12), .Z(n9) );
  CKBD1BWP U94 ( .I(n13), .Z(n8) );
  CKBD1BWP U95 ( .I(n14), .Z(n5) );
  CKBD1BWP U96 ( .I(n14), .Z(n3) );
  CKBD1BWP U97 ( .I(n14), .Z(n4) );
  CKBD1BWP U98 ( .I(n15), .Z(n1) );
  CKBD1BWP U99 ( .I(n15), .Z(n2) );
  CKBD1BWP U100 ( .I(n12), .Z(n11) );
  CKBD1BWP U101 ( .I(n172), .Z(n12) );
  CKBD1BWP U102 ( .I(n172), .Z(n13) );
  CKBD1BWP U103 ( .I(n172), .Z(n14) );
  CKBD1BWP U104 ( .I(n172), .Z(n15) );
  CKBD1BWP U105 ( .I(n42), .Z(n32) );
  CKBD1BWP U106 ( .I(n42), .Z(n33) );
  CKBD1BWP U107 ( .I(n42), .Z(n34) );
  CKBD1BWP U108 ( .I(n42), .Z(n35) );
  CKBD1BWP U109 ( .I(n42), .Z(n36) );
  CKBD1BWP U110 ( .I(n42), .Z(n37) );
  CKBD1BWP U111 ( .I(n42), .Z(n38) );
  CKBD1BWP U112 ( .I(n42), .Z(n39) );
  CKBD1BWP U113 ( .I(n42), .Z(n40) );
  CKBD1BWP U114 ( .I(n42), .Z(n41) );
  CKBD1BWP U115 ( .I(n28), .Z(n17) );
  CKBD1BWP U116 ( .I(n28), .Z(n18) );
  CKBD1BWP U117 ( .I(n28), .Z(n19) );
  CKBD1BWP U118 ( .I(n27), .Z(n20) );
  CKBD1BWP U119 ( .I(n27), .Z(n21) );
  CKBD1BWP U120 ( .I(n27), .Z(n22) );
  INVD1BWP U121 ( .I(\ML_int[7][127] ), .ZN(n43) );
  INVD1BWP U122 ( .I(\ML_int[7][126] ), .ZN(n44) );
  INVD1BWP U123 ( .I(\ML_int[7][125] ), .ZN(n45) );
  INVD1BWP U124 ( .I(\ML_int[7][124] ), .ZN(n46) );
  INVD1BWP U125 ( .I(\ML_int[7][123] ), .ZN(n47) );
  INVD1BWP U126 ( .I(\ML_int[7][122] ), .ZN(n48) );
  INVD1BWP U127 ( .I(\ML_int[7][121] ), .ZN(n49) );
  INVD1BWP U128 ( .I(\ML_int[7][120] ), .ZN(n50) );
  INVD1BWP U129 ( .I(\ML_int[7][119] ), .ZN(n51) );
  INVD1BWP U130 ( .I(\ML_int[7][118] ), .ZN(n52) );
  INVD1BWP U131 ( .I(\ML_int[7][117] ), .ZN(n53) );
  INVD1BWP U132 ( .I(\ML_int[7][116] ), .ZN(n54) );
  INVD1BWP U133 ( .I(\ML_int[7][115] ), .ZN(n55) );
  INVD1BWP U134 ( .I(\ML_int[7][114] ), .ZN(n56) );
  INVD1BWP U135 ( .I(\ML_int[7][113] ), .ZN(n57) );
  INVD1BWP U136 ( .I(\ML_int[7][112] ), .ZN(n58) );
  INVD1BWP U137 ( .I(\ML_int[7][111] ), .ZN(n59) );
  INVD1BWP U138 ( .I(\ML_int[7][110] ), .ZN(n60) );
  INVD1BWP U139 ( .I(\ML_int[7][109] ), .ZN(n61) );
  INVD1BWP U140 ( .I(\ML_int[7][108] ), .ZN(n62) );
  INVD1BWP U141 ( .I(\ML_int[7][107] ), .ZN(n63) );
  INVD1BWP U142 ( .I(\ML_int[7][106] ), .ZN(n64) );
  INVD1BWP U143 ( .I(\ML_int[7][105] ), .ZN(n65) );
  INVD1BWP U144 ( .I(\ML_int[7][104] ), .ZN(n66) );
  INVD1BWP U145 ( .I(\ML_int[7][103] ), .ZN(n67) );
  INVD1BWP U146 ( .I(\ML_int[7][102] ), .ZN(n68) );
  INVD1BWP U147 ( .I(\ML_int[7][101] ), .ZN(n69) );
  INVD1BWP U148 ( .I(\ML_int[7][100] ), .ZN(n70) );
  INVD1BWP U149 ( .I(\ML_int[7][99] ), .ZN(n71) );
  INVD1BWP U150 ( .I(\ML_int[7][98] ), .ZN(n72) );
  INVD1BWP U151 ( .I(\ML_int[7][97] ), .ZN(n73) );
  INVD1BWP U152 ( .I(\ML_int[7][96] ), .ZN(n74) );
  INVD1BWP U153 ( .I(\ML_int[7][95] ), .ZN(n75) );
  INVD1BWP U154 ( .I(\ML_int[7][94] ), .ZN(n76) );
  INVD1BWP U155 ( .I(\ML_int[7][93] ), .ZN(n77) );
  INVD1BWP U156 ( .I(\ML_int[7][92] ), .ZN(n78) );
  INVD1BWP U157 ( .I(\ML_int[7][91] ), .ZN(n79) );
  INVD1BWP U158 ( .I(\ML_int[7][90] ), .ZN(n80) );
  INVD1BWP U159 ( .I(\ML_int[7][89] ), .ZN(n81) );
  INVD1BWP U160 ( .I(\ML_int[7][88] ), .ZN(n82) );
  INVD1BWP U161 ( .I(\ML_int[7][87] ), .ZN(n83) );
  INVD1BWP U162 ( .I(\ML_int[7][86] ), .ZN(n84) );
  INVD1BWP U163 ( .I(\ML_int[7][85] ), .ZN(n85) );
  INVD1BWP U164 ( .I(\ML_int[7][84] ), .ZN(n86) );
  INVD1BWP U165 ( .I(\ML_int[7][83] ), .ZN(n87) );
  INVD1BWP U166 ( .I(\ML_int[7][82] ), .ZN(n88) );
  INVD1BWP U167 ( .I(\ML_int[7][81] ), .ZN(n89) );
  INVD1BWP U168 ( .I(\ML_int[7][80] ), .ZN(n90) );
  INVD1BWP U169 ( .I(\ML_int[7][79] ), .ZN(n91) );
  INVD1BWP U170 ( .I(\ML_int[7][78] ), .ZN(n92) );
  INVD1BWP U171 ( .I(\ML_int[7][77] ), .ZN(n93) );
  INVD1BWP U172 ( .I(\ML_int[7][76] ), .ZN(n94) );
  INVD1BWP U173 ( .I(\ML_int[7][75] ), .ZN(n95) );
  INVD1BWP U174 ( .I(\ML_int[7][74] ), .ZN(n96) );
  INVD1BWP U175 ( .I(\ML_int[7][73] ), .ZN(n97) );
  INVD1BWP U176 ( .I(\ML_int[7][72] ), .ZN(n98) );
  INVD1BWP U177 ( .I(\ML_int[7][71] ), .ZN(n99) );
  INVD1BWP U178 ( .I(\ML_int[7][70] ), .ZN(n100) );
  INVD1BWP U179 ( .I(\ML_int[7][69] ), .ZN(n101) );
  INVD1BWP U180 ( .I(\ML_int[7][68] ), .ZN(n102) );
  INVD1BWP U181 ( .I(\ML_int[7][67] ), .ZN(n103) );
  INVD1BWP U182 ( .I(\ML_int[7][66] ), .ZN(n104) );
  INVD1BWP U183 ( .I(\ML_int[7][65] ), .ZN(n105) );
  INVD1BWP U184 ( .I(\ML_int[7][64] ), .ZN(n106) );
  CKBD1BWP U185 ( .I(n30), .Z(n28) );
  CKBD1BWP U186 ( .I(n30), .Z(n27) );
  CKBD1BWP U187 ( .I(n26), .Z(n23) );
  CKBD1BWP U188 ( .I(n26), .Z(n24) );
  CKBD1BWP U189 ( .I(n29), .Z(n16) );
  CKBD1BWP U190 ( .I(n30), .Z(n29) );
  CKBD1BWP U191 ( .I(n26), .Z(n25) );
  INVD1BWP U192 ( .I(\temp_int_SH[7] ), .ZN(n42) );
  CKND1BWP U193 ( .I(\temp_int_SH[6] ), .ZN(n107) );
  AN2XD1BWP U194 ( .A1(\ML_int[6][63] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][127] ) );
  AN2XD1BWP U195 ( .A1(\ML_int[6][62] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][126] ) );
  AN2XD1BWP U196 ( .A1(\ML_int[6][61] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][125] ) );
  AN2XD1BWP U197 ( .A1(\ML_int[6][60] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][124] ) );
  AN2XD1BWP U198 ( .A1(\ML_int[6][59] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][123] ) );
  AN2XD1BWP U199 ( .A1(\ML_int[6][58] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][122] ) );
  AN2XD1BWP U200 ( .A1(\ML_int[6][57] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][121] ) );
  AN2XD1BWP U201 ( .A1(\ML_int[6][56] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][120] ) );
  AN2XD1BWP U202 ( .A1(\ML_int[6][55] ), .A2(\temp_int_SH[6] ), .Z(
        \ML_int[7][119] ) );
  CKBD1BWP U203 ( .I(n173), .Z(n30) );
  CKBD1BWP U204 ( .I(n31), .Z(n26) );
  CKBD1BWP U205 ( .I(n173), .Z(n31) );
  AN2XD1BWP U206 ( .A1(A[15]), .A2(\temp_int_SH[4] ), .Z(\ML_int[5][31] ) );
  AN2XD1BWP U207 ( .A1(A[14]), .A2(\temp_int_SH[4] ), .Z(\ML_int[5][30] ) );
  AN2XD1BWP U208 ( .A1(A[13]), .A2(\temp_int_SH[4] ), .Z(\ML_int[5][29] ) );
  AN2XD1BWP U209 ( .A1(A[12]), .A2(\temp_int_SH[4] ), .Z(\ML_int[5][28] ) );
  AN2XD1BWP U210 ( .A1(A[11]), .A2(\temp_int_SH[4] ), .Z(\ML_int[5][27] ) );
  AN2XD1BWP U211 ( .A1(A[10]), .A2(\temp_int_SH[4] ), .Z(\ML_int[5][26] ) );
  AN2XD1BWP U212 ( .A1(A[9]), .A2(\temp_int_SH[4] ), .Z(\ML_int[5][25] ) );
  AN2XD1BWP U213 ( .A1(A[8]), .A2(\temp_int_SH[4] ), .Z(\ML_int[5][24] ) );
  AN2XD1BWP U214 ( .A1(A[7]), .A2(\temp_int_SH[4] ), .Z(\ML_int[5][23] ) );
  AN2XD1BWP U215 ( .A1(A[6]), .A2(\temp_int_SH[4] ), .Z(\ML_int[5][22] ) );
  AN2XD1BWP U216 ( .A1(A[5]), .A2(\temp_int_SH[4] ), .Z(\ML_int[5][21] ) );
  AN2XD1BWP U217 ( .A1(A[4]), .A2(\temp_int_SH[4] ), .Z(\ML_int[5][20] ) );
  AN2XD1BWP U218 ( .A1(A[3]), .A2(\temp_int_SH[4] ), .Z(\ML_int[5][19] ) );
  AN2XD1BWP U219 ( .A1(A[2]), .A2(\temp_int_SH[4] ), .Z(\ML_int[5][18] ) );
  AN2XD1BWP U220 ( .A1(A[1]), .A2(\temp_int_SH[4] ), .Z(\ML_int[5][17] ) );
  AN2XD1BWP U221 ( .A1(\ML_int[4][0] ), .A2(\temp_int_SH[4] ), .Z(
        \ML_int[5][16] ) );
  NR2XD0BWP U222 ( .A1(n43), .A2(n32), .ZN(\ML_int[8][255] ) );
  NR2XD0BWP U223 ( .A1(n44), .A2(n32), .ZN(\ML_int[8][254] ) );
  NR2XD0BWP U224 ( .A1(n45), .A2(n32), .ZN(\ML_int[8][253] ) );
  NR2XD0BWP U225 ( .A1(n46), .A2(n32), .ZN(\ML_int[8][252] ) );
  NR2XD0BWP U226 ( .A1(n47), .A2(n32), .ZN(\ML_int[8][251] ) );
  NR2XD0BWP U227 ( .A1(n48), .A2(n32), .ZN(\ML_int[8][250] ) );
  NR2XD0BWP U228 ( .A1(n49), .A2(n32), .ZN(\ML_int[8][249] ) );
  NR2XD0BWP U229 ( .A1(n50), .A2(n32), .ZN(\ML_int[8][248] ) );
  NR2XD0BWP U230 ( .A1(n51), .A2(n32), .ZN(\ML_int[8][247] ) );
  NR2XD0BWP U231 ( .A1(n52), .A2(n32), .ZN(\ML_int[8][246] ) );
  NR2XD0BWP U232 ( .A1(n53), .A2(n32), .ZN(\ML_int[8][245] ) );
  NR2XD0BWP U233 ( .A1(n54), .A2(n32), .ZN(\ML_int[8][244] ) );
  NR2XD0BWP U234 ( .A1(n55), .A2(n32), .ZN(\ML_int[8][243] ) );
  NR2XD0BWP U235 ( .A1(n56), .A2(n33), .ZN(\ML_int[8][242] ) );
  NR2XD0BWP U236 ( .A1(n57), .A2(n33), .ZN(\ML_int[8][241] ) );
  NR2XD0BWP U237 ( .A1(n58), .A2(n33), .ZN(\ML_int[8][240] ) );
  NR2XD0BWP U238 ( .A1(n59), .A2(n33), .ZN(\ML_int[8][239] ) );
  NR2XD0BWP U239 ( .A1(n60), .A2(n33), .ZN(\ML_int[8][238] ) );
  NR2XD0BWP U240 ( .A1(n61), .A2(n33), .ZN(\ML_int[8][237] ) );
  NR2XD0BWP U241 ( .A1(n62), .A2(n33), .ZN(\ML_int[8][236] ) );
  NR2XD0BWP U242 ( .A1(n63), .A2(n33), .ZN(\ML_int[8][235] ) );
  NR2XD0BWP U243 ( .A1(n64), .A2(n33), .ZN(\ML_int[8][234] ) );
  NR2XD0BWP U244 ( .A1(n65), .A2(n33), .ZN(\ML_int[8][233] ) );
  NR2XD0BWP U245 ( .A1(n66), .A2(n33), .ZN(\ML_int[8][232] ) );
  NR2XD0BWP U246 ( .A1(n67), .A2(n33), .ZN(\ML_int[8][231] ) );
  NR2XD0BWP U247 ( .A1(n68), .A2(n33), .ZN(\ML_int[8][230] ) );
  NR2XD0BWP U248 ( .A1(n69), .A2(n34), .ZN(\ML_int[8][229] ) );
  NR2XD0BWP U249 ( .A1(n70), .A2(n34), .ZN(\ML_int[8][228] ) );
  NR2XD0BWP U250 ( .A1(n71), .A2(n34), .ZN(\ML_int[8][227] ) );
  NR2XD0BWP U251 ( .A1(n72), .A2(n34), .ZN(\ML_int[8][226] ) );
  NR2XD0BWP U252 ( .A1(n73), .A2(n34), .ZN(\ML_int[8][225] ) );
  NR2XD0BWP U253 ( .A1(n74), .A2(n34), .ZN(\ML_int[8][224] ) );
  NR2XD0BWP U254 ( .A1(n75), .A2(n34), .ZN(\ML_int[8][223] ) );
  NR2XD0BWP U255 ( .A1(n76), .A2(n34), .ZN(\ML_int[8][222] ) );
  NR2XD0BWP U256 ( .A1(n77), .A2(n34), .ZN(\ML_int[8][221] ) );
  NR2XD0BWP U257 ( .A1(n78), .A2(n34), .ZN(\ML_int[8][220] ) );
  NR2XD0BWP U258 ( .A1(n79), .A2(n34), .ZN(\ML_int[8][219] ) );
  NR2XD0BWP U259 ( .A1(n80), .A2(n34), .ZN(\ML_int[8][218] ) );
  NR2XD0BWP U260 ( .A1(n81), .A2(n34), .ZN(\ML_int[8][217] ) );
  NR2XD0BWP U261 ( .A1(n82), .A2(n35), .ZN(\ML_int[8][216] ) );
  NR2XD0BWP U262 ( .A1(n83), .A2(n35), .ZN(\ML_int[8][215] ) );
  NR2XD0BWP U263 ( .A1(n84), .A2(n35), .ZN(\ML_int[8][214] ) );
  NR2XD0BWP U264 ( .A1(n85), .A2(n35), .ZN(\ML_int[8][213] ) );
  NR2XD0BWP U265 ( .A1(n86), .A2(n35), .ZN(\ML_int[8][212] ) );
  NR2XD0BWP U266 ( .A1(n87), .A2(n35), .ZN(\ML_int[8][211] ) );
  NR2XD0BWP U267 ( .A1(n88), .A2(n35), .ZN(\ML_int[8][210] ) );
  NR2XD0BWP U268 ( .A1(n89), .A2(n35), .ZN(\ML_int[8][209] ) );
  NR2XD0BWP U269 ( .A1(n90), .A2(n35), .ZN(\ML_int[8][208] ) );
  NR2XD0BWP U270 ( .A1(n91), .A2(n35), .ZN(\ML_int[8][207] ) );
  NR2XD0BWP U271 ( .A1(n92), .A2(n35), .ZN(\ML_int[8][206] ) );
  NR2XD0BWP U272 ( .A1(n93), .A2(n35), .ZN(\ML_int[8][205] ) );
  NR2XD0BWP U273 ( .A1(n94), .A2(n35), .ZN(\ML_int[8][204] ) );
  NR2XD0BWP U274 ( .A1(n95), .A2(n36), .ZN(\ML_int[8][203] ) );
  NR2XD0BWP U275 ( .A1(n96), .A2(n36), .ZN(\ML_int[8][202] ) );
  NR2XD0BWP U276 ( .A1(n97), .A2(n36), .ZN(\ML_int[8][201] ) );
  NR2XD0BWP U277 ( .A1(n98), .A2(n36), .ZN(\ML_int[8][200] ) );
  NR2XD0BWP U278 ( .A1(n99), .A2(n36), .ZN(\ML_int[8][199] ) );
  NR2XD0BWP U279 ( .A1(n100), .A2(n36), .ZN(\ML_int[8][198] ) );
  NR2XD0BWP U280 ( .A1(n101), .A2(n36), .ZN(\ML_int[8][197] ) );
  NR2XD0BWP U281 ( .A1(n102), .A2(n36), .ZN(\ML_int[8][196] ) );
  NR2XD0BWP U282 ( .A1(n103), .A2(n36), .ZN(\ML_int[8][195] ) );
  NR2XD0BWP U283 ( .A1(n104), .A2(n36), .ZN(\ML_int[8][194] ) );
  NR2XD0BWP U284 ( .A1(n105), .A2(n36), .ZN(\ML_int[8][193] ) );
  NR2XD0BWP U285 ( .A1(n106), .A2(n36), .ZN(\ML_int[8][192] ) );
  NR2XD0BWP U286 ( .A1(n112), .A2(n36), .ZN(\ML_int[8][191] ) );
  NR2XD0BWP U287 ( .A1(n113), .A2(n37), .ZN(\ML_int[8][190] ) );
  NR2XD0BWP U288 ( .A1(n114), .A2(n37), .ZN(\ML_int[8][189] ) );
  NR2XD0BWP U289 ( .A1(n115), .A2(n37), .ZN(\ML_int[8][188] ) );
  NR2XD0BWP U290 ( .A1(n117), .A2(n37), .ZN(\ML_int[8][187] ) );
  NR2XD0BWP U291 ( .A1(n118), .A2(n37), .ZN(\ML_int[8][186] ) );
  NR2XD0BWP U292 ( .A1(n119), .A2(n37), .ZN(\ML_int[8][185] ) );
  NR2XD0BWP U293 ( .A1(n120), .A2(n37), .ZN(\ML_int[8][184] ) );
  NR2XD0BWP U294 ( .A1(n121), .A2(n37), .ZN(\ML_int[8][183] ) );
  NR2XD0BWP U295 ( .A1(n122), .A2(n37), .ZN(\ML_int[8][182] ) );
  NR2XD0BWP U296 ( .A1(n123), .A2(n37), .ZN(\ML_int[8][181] ) );
  NR2XD0BWP U297 ( .A1(n124), .A2(n37), .ZN(\ML_int[8][180] ) );
  NR2XD0BWP U298 ( .A1(n125), .A2(n37), .ZN(\ML_int[8][179] ) );
  NR2XD0BWP U299 ( .A1(n126), .A2(n37), .ZN(\ML_int[8][178] ) );
  NR2XD0BWP U300 ( .A1(n128), .A2(n38), .ZN(\ML_int[8][177] ) );
  NR2XD0BWP U301 ( .A1(n129), .A2(n38), .ZN(\ML_int[8][176] ) );
  NR2XD0BWP U302 ( .A1(n130), .A2(n38), .ZN(\ML_int[8][175] ) );
  NR2XD0BWP U303 ( .A1(n131), .A2(n38), .ZN(\ML_int[8][174] ) );
  NR2XD0BWP U304 ( .A1(n132), .A2(n38), .ZN(\ML_int[8][173] ) );
  NR2XD0BWP U305 ( .A1(n133), .A2(n38), .ZN(\ML_int[8][172] ) );
  NR2XD0BWP U306 ( .A1(n134), .A2(n38), .ZN(\ML_int[8][171] ) );
  NR2XD0BWP U307 ( .A1(n135), .A2(n38), .ZN(\ML_int[8][170] ) );
  NR2XD0BWP U308 ( .A1(n136), .A2(n38), .ZN(\ML_int[8][169] ) );
  NR2XD0BWP U309 ( .A1(n137), .A2(n38), .ZN(\ML_int[8][168] ) );
  NR2XD0BWP U310 ( .A1(n139), .A2(n38), .ZN(\ML_int[8][167] ) );
  NR2XD0BWP U311 ( .A1(n140), .A2(n38), .ZN(\ML_int[8][166] ) );
  NR2XD0BWP U312 ( .A1(n141), .A2(n38), .ZN(\ML_int[8][165] ) );
  NR2XD0BWP U313 ( .A1(n142), .A2(n39), .ZN(\ML_int[8][164] ) );
  NR2XD0BWP U314 ( .A1(n143), .A2(n39), .ZN(\ML_int[8][163] ) );
  NR2XD0BWP U315 ( .A1(n144), .A2(n39), .ZN(\ML_int[8][162] ) );
  NR2XD0BWP U316 ( .A1(n145), .A2(n39), .ZN(\ML_int[8][161] ) );
  NR2XD0BWP U317 ( .A1(n146), .A2(n39), .ZN(\ML_int[8][160] ) );
  NR2XD0BWP U318 ( .A1(n147), .A2(n39), .ZN(\ML_int[8][159] ) );
  NR2XD0BWP U319 ( .A1(n148), .A2(n39), .ZN(\ML_int[8][158] ) );
  NR2XD0BWP U320 ( .A1(n150), .A2(n39), .ZN(\ML_int[8][157] ) );
  NR2XD0BWP U321 ( .A1(n151), .A2(n39), .ZN(\ML_int[8][156] ) );
  NR2XD0BWP U322 ( .A1(n152), .A2(n39), .ZN(\ML_int[8][155] ) );
  NR2XD0BWP U323 ( .A1(n153), .A2(n39), .ZN(\ML_int[8][154] ) );
  NR2XD0BWP U324 ( .A1(n154), .A2(n39), .ZN(\ML_int[8][153] ) );
  NR2XD0BWP U325 ( .A1(n155), .A2(n39), .ZN(\ML_int[8][152] ) );
  NR2XD0BWP U326 ( .A1(n156), .A2(n40), .ZN(\ML_int[8][151] ) );
  NR2XD0BWP U327 ( .A1(n157), .A2(n40), .ZN(\ML_int[8][150] ) );
  NR2XD0BWP U328 ( .A1(n158), .A2(n40), .ZN(\ML_int[8][149] ) );
  NR2XD0BWP U329 ( .A1(n159), .A2(n40), .ZN(\ML_int[8][148] ) );
  NR2XD0BWP U330 ( .A1(n161), .A2(n40), .ZN(\ML_int[8][147] ) );
  NR2XD0BWP U331 ( .A1(n162), .A2(n40), .ZN(\ML_int[8][146] ) );
  NR2XD0BWP U332 ( .A1(n163), .A2(n40), .ZN(\ML_int[8][145] ) );
  NR2XD0BWP U333 ( .A1(n164), .A2(n40), .ZN(\ML_int[8][144] ) );
  NR2XD0BWP U334 ( .A1(n165), .A2(n40), .ZN(\ML_int[8][143] ) );
  NR2XD0BWP U335 ( .A1(n166), .A2(n40), .ZN(\ML_int[8][142] ) );
  NR2XD0BWP U336 ( .A1(n167), .A2(n40), .ZN(\ML_int[8][141] ) );
  NR2XD0BWP U337 ( .A1(n168), .A2(n40), .ZN(\ML_int[8][140] ) );
  NR2XD0BWP U338 ( .A1(n169), .A2(n40), .ZN(\ML_int[8][139] ) );
  NR2XD0BWP U339 ( .A1(n170), .A2(n41), .ZN(\ML_int[8][138] ) );
  NR2XD0BWP U340 ( .A1(n108), .A2(n41), .ZN(\ML_int[8][137] ) );
  NR2XD0BWP U341 ( .A1(n109), .A2(n41), .ZN(\ML_int[8][136] ) );
  NR2XD0BWP U342 ( .A1(n110), .A2(n41), .ZN(\ML_int[8][135] ) );
  NR2XD0BWP U343 ( .A1(n111), .A2(n41), .ZN(\ML_int[8][134] ) );
  NR2XD0BWP U344 ( .A1(n116), .A2(n41), .ZN(\ML_int[8][133] ) );
  NR2XD0BWP U345 ( .A1(n127), .A2(n41), .ZN(\ML_int[8][132] ) );
  NR2XD0BWP U346 ( .A1(n138), .A2(n41), .ZN(\ML_int[8][131] ) );
  NR2XD0BWP U347 ( .A1(n149), .A2(n41), .ZN(\ML_int[8][130] ) );
  NR2XD0BWP U348 ( .A1(n160), .A2(n41), .ZN(\ML_int[8][129] ) );
  NR2XD0BWP U349 ( .A1(n171), .A2(n41), .ZN(\ML_int[8][128] ) );
  NR2D0BWP U350 ( .A1(n1), .A2(n108), .ZN(\ML_int[10][9] ) );
  CKND2D0BWP U351 ( .A1(\ML_int[6][9] ), .A2(n107), .ZN(n108) );
  INR2D0BWP U352 ( .A1(\ML_int[5][9] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][9] ) );
  INR2D0BWP U353 ( .A1(A[9]), .B1(\temp_int_SH[4] ), .ZN(\ML_int[5][9] ) );
  INR2D0BWP U354 ( .A1(\ML_int[7][99] ), .B1(n11), .ZN(\ML_int[10][99] ) );
  INR2D0BWP U355 ( .A1(\ML_int[7][98] ), .B1(n11), .ZN(\ML_int[10][98] ) );
  INR2D0BWP U356 ( .A1(\ML_int[7][97] ), .B1(n10), .ZN(\ML_int[10][97] ) );
  INR2D0BWP U357 ( .A1(\ML_int[7][96] ), .B1(n10), .ZN(\ML_int[10][96] ) );
  INR2D0BWP U358 ( .A1(\ML_int[7][95] ), .B1(n10), .ZN(\ML_int[10][95] ) );
  INR2D0BWP U359 ( .A1(\ML_int[7][94] ), .B1(n10), .ZN(\ML_int[10][94] ) );
  INR2D0BWP U360 ( .A1(\ML_int[7][93] ), .B1(n10), .ZN(\ML_int[10][93] ) );
  INR2D0BWP U361 ( .A1(\ML_int[7][92] ), .B1(n10), .ZN(\ML_int[10][92] ) );
  INR2D0BWP U362 ( .A1(\ML_int[7][91] ), .B1(n10), .ZN(\ML_int[10][91] ) );
  INR2D0BWP U363 ( .A1(\ML_int[7][90] ), .B1(n10), .ZN(\ML_int[10][90] ) );
  NR2D0BWP U364 ( .A1(n1), .A2(n109), .ZN(\ML_int[10][8] ) );
  CKND2D0BWP U365 ( .A1(\ML_int[6][8] ), .A2(n107), .ZN(n109) );
  INR2D0BWP U366 ( .A1(\ML_int[5][8] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][8] ) );
  INR2D0BWP U367 ( .A1(A[8]), .B1(\temp_int_SH[4] ), .ZN(\ML_int[5][8] ) );
  INR2D0BWP U368 ( .A1(\ML_int[7][89] ), .B1(n10), .ZN(\ML_int[10][89] ) );
  INR2D0BWP U369 ( .A1(\ML_int[7][88] ), .B1(n10), .ZN(\ML_int[10][88] ) );
  INR2D0BWP U370 ( .A1(\ML_int[7][87] ), .B1(n10), .ZN(\ML_int[10][87] ) );
  INR2D0BWP U371 ( .A1(\ML_int[7][86] ), .B1(n10), .ZN(\ML_int[10][86] ) );
  INR2D0BWP U372 ( .A1(\ML_int[7][85] ), .B1(n9), .ZN(\ML_int[10][85] ) );
  INR2D0BWP U373 ( .A1(\ML_int[7][84] ), .B1(n9), .ZN(\ML_int[10][84] ) );
  INR2D0BWP U374 ( .A1(\ML_int[7][83] ), .B1(n9), .ZN(\ML_int[10][83] ) );
  INR2D0BWP U375 ( .A1(\ML_int[7][82] ), .B1(n9), .ZN(\ML_int[10][82] ) );
  INR2D0BWP U376 ( .A1(\ML_int[7][81] ), .B1(n9), .ZN(\ML_int[10][81] ) );
  INR2D0BWP U377 ( .A1(\ML_int[7][80] ), .B1(n9), .ZN(\ML_int[10][80] ) );
  NR2D0BWP U378 ( .A1(n1), .A2(n110), .ZN(\ML_int[10][7] ) );
  CKND2D0BWP U379 ( .A1(\ML_int[6][7] ), .A2(n107), .ZN(n110) );
  INR2D0BWP U380 ( .A1(\ML_int[5][7] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][7] ) );
  INR2D0BWP U381 ( .A1(A[7]), .B1(\temp_int_SH[4] ), .ZN(\ML_int[5][7] ) );
  INR2D0BWP U382 ( .A1(\ML_int[7][79] ), .B1(n9), .ZN(\ML_int[10][79] ) );
  INR2D0BWP U383 ( .A1(\ML_int[7][78] ), .B1(n9), .ZN(\ML_int[10][78] ) );
  INR2D0BWP U384 ( .A1(\ML_int[7][77] ), .B1(n9), .ZN(\ML_int[10][77] ) );
  INR2D0BWP U385 ( .A1(\ML_int[7][76] ), .B1(n9), .ZN(\ML_int[10][76] ) );
  INR2D0BWP U386 ( .A1(\ML_int[7][75] ), .B1(n9), .ZN(\ML_int[10][75] ) );
  INR2D0BWP U387 ( .A1(\ML_int[7][74] ), .B1(n9), .ZN(\ML_int[10][74] ) );
  INR2D0BWP U388 ( .A1(\ML_int[7][73] ), .B1(n8), .ZN(\ML_int[10][73] ) );
  INR2D0BWP U389 ( .A1(\ML_int[7][72] ), .B1(n8), .ZN(\ML_int[10][72] ) );
  INR2D0BWP U390 ( .A1(\ML_int[7][71] ), .B1(n8), .ZN(\ML_int[10][71] ) );
  INR2D0BWP U391 ( .A1(\ML_int[7][70] ), .B1(n8), .ZN(\ML_int[10][70] ) );
  NR2D0BWP U392 ( .A1(n1), .A2(n111), .ZN(\ML_int[10][6] ) );
  CKND2D0BWP U393 ( .A1(\ML_int[6][6] ), .A2(n107), .ZN(n111) );
  INR2D0BWP U394 ( .A1(\ML_int[5][6] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][6] ) );
  INR2D0BWP U395 ( .A1(A[6]), .B1(\temp_int_SH[4] ), .ZN(\ML_int[5][6] ) );
  INR2D0BWP U396 ( .A1(\ML_int[7][69] ), .B1(n8), .ZN(\ML_int[10][69] ) );
  INR2D0BWP U397 ( .A1(\ML_int[7][68] ), .B1(n8), .ZN(\ML_int[10][68] ) );
  INR2D0BWP U398 ( .A1(\ML_int[7][67] ), .B1(n8), .ZN(\ML_int[10][67] ) );
  INR2D0BWP U399 ( .A1(\ML_int[7][66] ), .B1(n8), .ZN(\ML_int[10][66] ) );
  INR2D0BWP U400 ( .A1(\ML_int[7][65] ), .B1(n8), .ZN(\ML_int[10][65] ) );
  INR2D0BWP U401 ( .A1(\ML_int[7][64] ), .B1(n8), .ZN(\ML_int[10][64] ) );
  NR2D0BWP U402 ( .A1(n1), .A2(n112), .ZN(\ML_int[10][63] ) );
  CKND2D0BWP U403 ( .A1(\ML_int[6][63] ), .A2(n107), .ZN(n112) );
  NR2D0BWP U404 ( .A1(n1), .A2(n113), .ZN(\ML_int[10][62] ) );
  CKND2D0BWP U405 ( .A1(\ML_int[6][62] ), .A2(n107), .ZN(n113) );
  NR2D0BWP U406 ( .A1(n1), .A2(n114), .ZN(\ML_int[10][61] ) );
  CKND2D0BWP U407 ( .A1(\ML_int[6][61] ), .A2(n107), .ZN(n114) );
  NR2D0BWP U408 ( .A1(n1), .A2(n115), .ZN(\ML_int[10][60] ) );
  CKND2D0BWP U409 ( .A1(\ML_int[6][60] ), .A2(n107), .ZN(n115) );
  NR2D0BWP U410 ( .A1(n1), .A2(n116), .ZN(\ML_int[10][5] ) );
  CKND2D0BWP U411 ( .A1(\ML_int[6][5] ), .A2(n107), .ZN(n116) );
  INR2D0BWP U412 ( .A1(\ML_int[5][5] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][5] ) );
  INR2D0BWP U413 ( .A1(A[5]), .B1(\temp_int_SH[4] ), .ZN(\ML_int[5][5] ) );
  NR2D0BWP U414 ( .A1(n1), .A2(n117), .ZN(\ML_int[10][59] ) );
  CKND2D0BWP U415 ( .A1(\ML_int[6][59] ), .A2(n107), .ZN(n117) );
  NR2D0BWP U416 ( .A1(n1), .A2(n118), .ZN(\ML_int[10][58] ) );
  CKND2D0BWP U417 ( .A1(\ML_int[6][58] ), .A2(n107), .ZN(n118) );
  NR2D0BWP U418 ( .A1(n1), .A2(n119), .ZN(\ML_int[10][57] ) );
  CKND2D0BWP U419 ( .A1(\ML_int[6][57] ), .A2(n107), .ZN(n119) );
  NR2D0BWP U420 ( .A1(n2), .A2(n120), .ZN(\ML_int[10][56] ) );
  CKND2D0BWP U421 ( .A1(\ML_int[6][56] ), .A2(n107), .ZN(n120) );
  NR2D0BWP U422 ( .A1(n2), .A2(n121), .ZN(\ML_int[10][55] ) );
  CKND2D0BWP U423 ( .A1(\ML_int[6][55] ), .A2(n107), .ZN(n121) );
  NR2D0BWP U424 ( .A1(n2), .A2(n122), .ZN(\ML_int[10][54] ) );
  CKND2D0BWP U425 ( .A1(\ML_int[6][54] ), .A2(n107), .ZN(n122) );
  NR2D0BWP U426 ( .A1(n2), .A2(n123), .ZN(\ML_int[10][53] ) );
  CKND2D0BWP U427 ( .A1(\ML_int[6][53] ), .A2(n107), .ZN(n123) );
  NR2D0BWP U428 ( .A1(n2), .A2(n124), .ZN(\ML_int[10][52] ) );
  CKND2D0BWP U429 ( .A1(\ML_int[6][52] ), .A2(n107), .ZN(n124) );
  NR2D0BWP U430 ( .A1(n2), .A2(n125), .ZN(\ML_int[10][51] ) );
  CKND2D0BWP U431 ( .A1(\ML_int[6][51] ), .A2(n107), .ZN(n125) );
  NR2D0BWP U432 ( .A1(n2), .A2(n126), .ZN(\ML_int[10][50] ) );
  CKND2D0BWP U433 ( .A1(\ML_int[6][50] ), .A2(n107), .ZN(n126) );
  NR2D0BWP U434 ( .A1(n2), .A2(n127), .ZN(\ML_int[10][4] ) );
  CKND2D0BWP U435 ( .A1(\ML_int[6][4] ), .A2(n107), .ZN(n127) );
  INR2D0BWP U436 ( .A1(\ML_int[5][4] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][4] ) );
  INR2D0BWP U437 ( .A1(A[4]), .B1(\temp_int_SH[4] ), .ZN(\ML_int[5][4] ) );
  NR2D0BWP U438 ( .A1(n2), .A2(n128), .ZN(\ML_int[10][49] ) );
  CKND2D0BWP U439 ( .A1(\ML_int[6][49] ), .A2(n107), .ZN(n128) );
  NR2D0BWP U440 ( .A1(n2), .A2(n129), .ZN(\ML_int[10][48] ) );
  CKND2D0BWP U441 ( .A1(\ML_int[6][48] ), .A2(n107), .ZN(n129) );
  NR2D0BWP U442 ( .A1(n2), .A2(n130), .ZN(\ML_int[10][47] ) );
  CKND2D0BWP U443 ( .A1(\ML_int[6][47] ), .A2(n107), .ZN(n130) );
  NR2D0BWP U444 ( .A1(n2), .A2(n131), .ZN(\ML_int[10][46] ) );
  CKND2D0BWP U445 ( .A1(\ML_int[6][46] ), .A2(n107), .ZN(n131) );
  NR2D0BWP U446 ( .A1(n3), .A2(n132), .ZN(\ML_int[10][45] ) );
  CKND2D0BWP U447 ( .A1(\ML_int[6][45] ), .A2(n107), .ZN(n132) );
  NR2D0BWP U448 ( .A1(n3), .A2(n133), .ZN(\ML_int[10][44] ) );
  CKND2D0BWP U449 ( .A1(\ML_int[6][44] ), .A2(n107), .ZN(n133) );
  NR2D0BWP U450 ( .A1(n3), .A2(n134), .ZN(\ML_int[10][43] ) );
  CKND2D0BWP U451 ( .A1(\ML_int[6][43] ), .A2(n107), .ZN(n134) );
  NR2D0BWP U452 ( .A1(n3), .A2(n135), .ZN(\ML_int[10][42] ) );
  CKND2D0BWP U453 ( .A1(\ML_int[6][42] ), .A2(n107), .ZN(n135) );
  NR2D0BWP U454 ( .A1(n3), .A2(n136), .ZN(\ML_int[10][41] ) );
  CKND2D0BWP U455 ( .A1(\ML_int[6][41] ), .A2(n107), .ZN(n136) );
  NR2D0BWP U456 ( .A1(n3), .A2(n137), .ZN(\ML_int[10][40] ) );
  CKND2D0BWP U457 ( .A1(\ML_int[6][40] ), .A2(n107), .ZN(n137) );
  NR2D0BWP U458 ( .A1(n3), .A2(n138), .ZN(\ML_int[10][3] ) );
  CKND2D0BWP U459 ( .A1(\ML_int[6][3] ), .A2(n107), .ZN(n138) );
  INR2D0BWP U460 ( .A1(\ML_int[5][3] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][3] ) );
  INR2D0BWP U461 ( .A1(A[3]), .B1(\temp_int_SH[4] ), .ZN(\ML_int[5][3] ) );
  NR2D0BWP U462 ( .A1(n3), .A2(n139), .ZN(\ML_int[10][39] ) );
  CKND2D0BWP U463 ( .A1(\ML_int[6][39] ), .A2(n107), .ZN(n139) );
  NR2D0BWP U464 ( .A1(n3), .A2(n140), .ZN(\ML_int[10][38] ) );
  CKND2D0BWP U465 ( .A1(\ML_int[6][38] ), .A2(n107), .ZN(n140) );
  NR2D0BWP U466 ( .A1(n3), .A2(n141), .ZN(\ML_int[10][37] ) );
  CKND2D0BWP U467 ( .A1(\ML_int[6][37] ), .A2(n107), .ZN(n141) );
  NR2D0BWP U468 ( .A1(n3), .A2(n142), .ZN(\ML_int[10][36] ) );
  CKND2D0BWP U469 ( .A1(\ML_int[6][36] ), .A2(n107), .ZN(n142) );
  NR2D0BWP U470 ( .A1(n3), .A2(n143), .ZN(\ML_int[10][35] ) );
  CKND2D0BWP U471 ( .A1(\ML_int[6][35] ), .A2(n107), .ZN(n143) );
  NR2D0BWP U472 ( .A1(n4), .A2(n144), .ZN(\ML_int[10][34] ) );
  CKND2D0BWP U473 ( .A1(\ML_int[6][34] ), .A2(n107), .ZN(n144) );
  NR2D0BWP U474 ( .A1(n4), .A2(n145), .ZN(\ML_int[10][33] ) );
  CKND2D0BWP U475 ( .A1(\ML_int[6][33] ), .A2(n107), .ZN(n145) );
  NR2D0BWP U476 ( .A1(n4), .A2(n146), .ZN(\ML_int[10][32] ) );
  CKND2D0BWP U477 ( .A1(\ML_int[6][32] ), .A2(n107), .ZN(n146) );
  NR2D0BWP U478 ( .A1(n4), .A2(n147), .ZN(\ML_int[10][31] ) );
  CKND2D0BWP U479 ( .A1(\ML_int[6][31] ), .A2(n107), .ZN(n147) );
  INR2D0BWP U480 ( .A1(\ML_int[5][31] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][31] ) );
  NR2D0BWP U481 ( .A1(n4), .A2(n148), .ZN(\ML_int[10][30] ) );
  CKND2D0BWP U482 ( .A1(\ML_int[6][30] ), .A2(n107), .ZN(n148) );
  INR2D0BWP U483 ( .A1(\ML_int[5][30] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][30] ) );
  NR2D0BWP U484 ( .A1(n4), .A2(n149), .ZN(\ML_int[10][2] ) );
  CKND2D0BWP U485 ( .A1(\ML_int[6][2] ), .A2(n107), .ZN(n149) );
  INR2D0BWP U486 ( .A1(\ML_int[5][2] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][2] ) );
  INR2D0BWP U487 ( .A1(A[2]), .B1(\temp_int_SH[4] ), .ZN(\ML_int[5][2] ) );
  NR2D0BWP U488 ( .A1(n4), .A2(n150), .ZN(\ML_int[10][29] ) );
  CKND2D0BWP U489 ( .A1(\ML_int[6][29] ), .A2(n107), .ZN(n150) );
  INR2D0BWP U490 ( .A1(\ML_int[5][29] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][29] ) );
  NR2D0BWP U491 ( .A1(n4), .A2(n151), .ZN(\ML_int[10][28] ) );
  CKND2D0BWP U492 ( .A1(\ML_int[6][28] ), .A2(n107), .ZN(n151) );
  INR2D0BWP U493 ( .A1(\ML_int[5][28] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][28] ) );
  NR2D0BWP U494 ( .A1(n4), .A2(n152), .ZN(\ML_int[10][27] ) );
  CKND2D0BWP U495 ( .A1(\ML_int[6][27] ), .A2(n107), .ZN(n152) );
  INR2D0BWP U496 ( .A1(\ML_int[5][27] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][27] ) );
  NR2D0BWP U497 ( .A1(n4), .A2(n153), .ZN(\ML_int[10][26] ) );
  CKND2D0BWP U498 ( .A1(\ML_int[6][26] ), .A2(n107), .ZN(n153) );
  INR2D0BWP U499 ( .A1(\ML_int[5][26] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][26] ) );
  NR2D0BWP U500 ( .A1(n4), .A2(n154), .ZN(\ML_int[10][25] ) );
  CKND2D0BWP U501 ( .A1(\ML_int[6][25] ), .A2(n107), .ZN(n154) );
  INR2D0BWP U502 ( .A1(\ML_int[5][25] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][25] ) );
  AN2D0BWP U503 ( .A1(\ML_int[8][255] ), .A2(n16), .Z(\ML_int[10][255] ) );
  AN2D0BWP U504 ( .A1(\ML_int[8][254] ), .A2(n16), .Z(\ML_int[10][254] ) );
  AN2D0BWP U505 ( .A1(\ML_int[8][253] ), .A2(n16), .Z(\ML_int[10][253] ) );
  AN2D0BWP U506 ( .A1(\ML_int[8][252] ), .A2(n16), .Z(\ML_int[10][252] ) );
  AN2D0BWP U507 ( .A1(\ML_int[8][251] ), .A2(n16), .Z(\ML_int[10][251] ) );
  AN2D0BWP U508 ( .A1(\ML_int[8][250] ), .A2(n16), .Z(\ML_int[10][250] ) );
  NR2D0BWP U509 ( .A1(n5), .A2(n155), .ZN(\ML_int[10][24] ) );
  CKND2D0BWP U510 ( .A1(\ML_int[6][24] ), .A2(n107), .ZN(n155) );
  INR2D0BWP U511 ( .A1(\ML_int[5][24] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][24] ) );
  AN2D0BWP U512 ( .A1(\ML_int[8][249] ), .A2(n16), .Z(\ML_int[10][249] ) );
  AN2D0BWP U513 ( .A1(\ML_int[8][248] ), .A2(n16), .Z(\ML_int[10][248] ) );
  AN2D0BWP U514 ( .A1(\ML_int[8][247] ), .A2(n16), .Z(\ML_int[10][247] ) );
  AN2D0BWP U515 ( .A1(\ML_int[8][246] ), .A2(n16), .Z(\ML_int[10][246] ) );
  AN2D0BWP U516 ( .A1(\ML_int[8][245] ), .A2(n16), .Z(\ML_int[10][245] ) );
  AN2D0BWP U517 ( .A1(\ML_int[8][244] ), .A2(n16), .Z(\ML_int[10][244] ) );
  AN2D0BWP U518 ( .A1(\ML_int[8][243] ), .A2(n16), .Z(\ML_int[10][243] ) );
  AN2D0BWP U519 ( .A1(\ML_int[8][242] ), .A2(n17), .Z(\ML_int[10][242] ) );
  AN2D0BWP U520 ( .A1(\ML_int[8][241] ), .A2(n17), .Z(\ML_int[10][241] ) );
  AN2D0BWP U521 ( .A1(\ML_int[8][240] ), .A2(n17), .Z(\ML_int[10][240] ) );
  NR2D0BWP U522 ( .A1(n5), .A2(n156), .ZN(\ML_int[10][23] ) );
  CKND2D0BWP U523 ( .A1(\ML_int[6][23] ), .A2(n107), .ZN(n156) );
  INR2D0BWP U524 ( .A1(\ML_int[5][23] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][23] ) );
  AN2D0BWP U525 ( .A1(\ML_int[8][239] ), .A2(n17), .Z(\ML_int[10][239] ) );
  AN2D0BWP U526 ( .A1(\ML_int[8][238] ), .A2(n17), .Z(\ML_int[10][238] ) );
  AN2D0BWP U527 ( .A1(\ML_int[8][237] ), .A2(n17), .Z(\ML_int[10][237] ) );
  AN2D0BWP U528 ( .A1(\ML_int[8][236] ), .A2(n17), .Z(\ML_int[10][236] ) );
  AN2D0BWP U529 ( .A1(\ML_int[8][235] ), .A2(n17), .Z(\ML_int[10][235] ) );
  AN2D0BWP U530 ( .A1(\ML_int[8][234] ), .A2(n17), .Z(\ML_int[10][234] ) );
  AN2D0BWP U531 ( .A1(\ML_int[8][233] ), .A2(n17), .Z(\ML_int[10][233] ) );
  AN2D0BWP U532 ( .A1(\ML_int[8][232] ), .A2(n17), .Z(\ML_int[10][232] ) );
  AN2D0BWP U533 ( .A1(\ML_int[8][231] ), .A2(n17), .Z(\ML_int[10][231] ) );
  AN2D0BWP U534 ( .A1(\ML_int[8][230] ), .A2(n17), .Z(\ML_int[10][230] ) );
  NR2D0BWP U535 ( .A1(n5), .A2(n157), .ZN(\ML_int[10][22] ) );
  CKND2D0BWP U536 ( .A1(\ML_int[6][22] ), .A2(n107), .ZN(n157) );
  INR2D0BWP U537 ( .A1(\ML_int[5][22] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][22] ) );
  AN2D0BWP U538 ( .A1(\ML_int[8][229] ), .A2(n18), .Z(\ML_int[10][229] ) );
  AN2D0BWP U539 ( .A1(\ML_int[8][228] ), .A2(n18), .Z(\ML_int[10][228] ) );
  AN2D0BWP U540 ( .A1(\ML_int[8][227] ), .A2(n18), .Z(\ML_int[10][227] ) );
  AN2D0BWP U541 ( .A1(\ML_int[8][226] ), .A2(n18), .Z(\ML_int[10][226] ) );
  AN2D0BWP U542 ( .A1(\ML_int[8][225] ), .A2(n18), .Z(\ML_int[10][225] ) );
  AN2D0BWP U543 ( .A1(\ML_int[8][224] ), .A2(n18), .Z(\ML_int[10][224] ) );
  AN2D0BWP U544 ( .A1(\ML_int[8][223] ), .A2(n18), .Z(\ML_int[10][223] ) );
  AN2D0BWP U545 ( .A1(\ML_int[8][222] ), .A2(n18), .Z(\ML_int[10][222] ) );
  AN2D0BWP U546 ( .A1(\ML_int[8][221] ), .A2(n18), .Z(\ML_int[10][221] ) );
  AN2D0BWP U547 ( .A1(\ML_int[8][220] ), .A2(n18), .Z(\ML_int[10][220] ) );
  NR2D0BWP U548 ( .A1(n5), .A2(n158), .ZN(\ML_int[10][21] ) );
  CKND2D0BWP U549 ( .A1(\ML_int[6][21] ), .A2(n107), .ZN(n158) );
  INR2D0BWP U550 ( .A1(\ML_int[5][21] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][21] ) );
  AN2D0BWP U551 ( .A1(\ML_int[8][219] ), .A2(n18), .Z(\ML_int[10][219] ) );
  AN2D0BWP U552 ( .A1(\ML_int[8][218] ), .A2(n18), .Z(\ML_int[10][218] ) );
  AN2D0BWP U553 ( .A1(\ML_int[8][217] ), .A2(n18), .Z(\ML_int[10][217] ) );
  AN2D0BWP U554 ( .A1(\ML_int[8][216] ), .A2(n19), .Z(\ML_int[10][216] ) );
  AN2D0BWP U555 ( .A1(\ML_int[8][215] ), .A2(n19), .Z(\ML_int[10][215] ) );
  AN2D0BWP U556 ( .A1(\ML_int[8][214] ), .A2(n19), .Z(\ML_int[10][214] ) );
  AN2D0BWP U557 ( .A1(\ML_int[8][213] ), .A2(n19), .Z(\ML_int[10][213] ) );
  AN2D0BWP U558 ( .A1(\ML_int[8][212] ), .A2(n19), .Z(\ML_int[10][212] ) );
  AN2D0BWP U559 ( .A1(\ML_int[8][211] ), .A2(n19), .Z(\ML_int[10][211] ) );
  AN2D0BWP U560 ( .A1(\ML_int[8][210] ), .A2(n19), .Z(\ML_int[10][210] ) );
  NR2D0BWP U561 ( .A1(n5), .A2(n159), .ZN(\ML_int[10][20] ) );
  CKND2D0BWP U562 ( .A1(\ML_int[6][20] ), .A2(n107), .ZN(n159) );
  INR2D0BWP U563 ( .A1(\ML_int[5][20] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][20] ) );
  AN2D0BWP U564 ( .A1(\ML_int[8][209] ), .A2(n19), .Z(\ML_int[10][209] ) );
  AN2D0BWP U565 ( .A1(\ML_int[8][208] ), .A2(n19), .Z(\ML_int[10][208] ) );
  AN2D0BWP U566 ( .A1(\ML_int[8][207] ), .A2(n19), .Z(\ML_int[10][207] ) );
  AN2D0BWP U567 ( .A1(\ML_int[8][206] ), .A2(n19), .Z(\ML_int[10][206] ) );
  AN2D0BWP U568 ( .A1(\ML_int[8][205] ), .A2(n19), .Z(\ML_int[10][205] ) );
  AN2D0BWP U569 ( .A1(\ML_int[8][204] ), .A2(n19), .Z(\ML_int[10][204] ) );
  AN2D0BWP U570 ( .A1(\ML_int[8][203] ), .A2(n20), .Z(\ML_int[10][203] ) );
  AN2D0BWP U571 ( .A1(\ML_int[8][202] ), .A2(n20), .Z(\ML_int[10][202] ) );
  AN2D0BWP U572 ( .A1(\ML_int[8][201] ), .A2(n20), .Z(\ML_int[10][201] ) );
  AN2D0BWP U573 ( .A1(\ML_int[8][200] ), .A2(n20), .Z(\ML_int[10][200] ) );
  NR2D0BWP U574 ( .A1(n5), .A2(n160), .ZN(\ML_int[10][1] ) );
  CKND2D0BWP U575 ( .A1(\ML_int[6][1] ), .A2(n107), .ZN(n160) );
  INR2D0BWP U576 ( .A1(\ML_int[5][1] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][1] ) );
  INR2D0BWP U577 ( .A1(A[1]), .B1(\temp_int_SH[4] ), .ZN(\ML_int[5][1] ) );
  NR2D0BWP U578 ( .A1(n5), .A2(n161), .ZN(\ML_int[10][19] ) );
  CKND2D0BWP U579 ( .A1(\ML_int[6][19] ), .A2(n107), .ZN(n161) );
  INR2D0BWP U580 ( .A1(\ML_int[5][19] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][19] ) );
  AN2D0BWP U581 ( .A1(\ML_int[8][199] ), .A2(n20), .Z(\ML_int[10][199] ) );
  AN2D0BWP U582 ( .A1(\ML_int[8][198] ), .A2(n20), .Z(\ML_int[10][198] ) );
  AN2D0BWP U583 ( .A1(\ML_int[8][197] ), .A2(n20), .Z(\ML_int[10][197] ) );
  AN2D0BWP U584 ( .A1(\ML_int[8][196] ), .A2(n20), .Z(\ML_int[10][196] ) );
  AN2D0BWP U585 ( .A1(\ML_int[8][195] ), .A2(n20), .Z(\ML_int[10][195] ) );
  AN2D0BWP U586 ( .A1(\ML_int[8][194] ), .A2(n20), .Z(\ML_int[10][194] ) );
  AN2D0BWP U587 ( .A1(\ML_int[8][193] ), .A2(n20), .Z(\ML_int[10][193] ) );
  AN2D0BWP U588 ( .A1(\ML_int[8][192] ), .A2(n20), .Z(\ML_int[10][192] ) );
  AN2D0BWP U589 ( .A1(\ML_int[8][191] ), .A2(n20), .Z(\ML_int[10][191] ) );
  AN2D0BWP U590 ( .A1(\ML_int[8][190] ), .A2(n21), .Z(\ML_int[10][190] ) );
  NR2D0BWP U591 ( .A1(n5), .A2(n162), .ZN(\ML_int[10][18] ) );
  CKND2D0BWP U592 ( .A1(\ML_int[6][18] ), .A2(n107), .ZN(n162) );
  INR2D0BWP U593 ( .A1(\ML_int[5][18] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][18] ) );
  AN2D0BWP U594 ( .A1(\ML_int[8][189] ), .A2(n21), .Z(\ML_int[10][189] ) );
  AN2D0BWP U595 ( .A1(\ML_int[8][188] ), .A2(n21), .Z(\ML_int[10][188] ) );
  AN2D0BWP U596 ( .A1(\ML_int[8][187] ), .A2(n21), .Z(\ML_int[10][187] ) );
  AN2D0BWP U597 ( .A1(\ML_int[8][186] ), .A2(n21), .Z(\ML_int[10][186] ) );
  AN2D0BWP U598 ( .A1(\ML_int[8][185] ), .A2(n21), .Z(\ML_int[10][185] ) );
  AN2D0BWP U599 ( .A1(\ML_int[8][184] ), .A2(n21), .Z(\ML_int[10][184] ) );
  AN2D0BWP U600 ( .A1(\ML_int[8][183] ), .A2(n21), .Z(\ML_int[10][183] ) );
  AN2D0BWP U601 ( .A1(\ML_int[8][182] ), .A2(n21), .Z(\ML_int[10][182] ) );
  AN2D0BWP U602 ( .A1(\ML_int[8][181] ), .A2(n21), .Z(\ML_int[10][181] ) );
  AN2D0BWP U603 ( .A1(\ML_int[8][180] ), .A2(n21), .Z(\ML_int[10][180] ) );
  NR2D0BWP U604 ( .A1(n5), .A2(n163), .ZN(\ML_int[10][17] ) );
  CKND2D0BWP U605 ( .A1(\ML_int[6][17] ), .A2(n107), .ZN(n163) );
  INR2D0BWP U606 ( .A1(\ML_int[5][17] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][17] ) );
  AN2D0BWP U607 ( .A1(\ML_int[8][179] ), .A2(n21), .Z(\ML_int[10][179] ) );
  AN2D0BWP U608 ( .A1(\ML_int[8][178] ), .A2(n21), .Z(\ML_int[10][178] ) );
  AN2D0BWP U609 ( .A1(\ML_int[8][177] ), .A2(n22), .Z(\ML_int[10][177] ) );
  AN2D0BWP U610 ( .A1(\ML_int[8][176] ), .A2(n22), .Z(\ML_int[10][176] ) );
  AN2D0BWP U611 ( .A1(\ML_int[8][175] ), .A2(n22), .Z(\ML_int[10][175] ) );
  AN2D0BWP U612 ( .A1(\ML_int[8][174] ), .A2(n22), .Z(\ML_int[10][174] ) );
  AN2D0BWP U613 ( .A1(\ML_int[8][173] ), .A2(n22), .Z(\ML_int[10][173] ) );
  AN2D0BWP U614 ( .A1(\ML_int[8][172] ), .A2(n22), .Z(\ML_int[10][172] ) );
  AN2D0BWP U615 ( .A1(\ML_int[8][171] ), .A2(n22), .Z(\ML_int[10][171] ) );
  AN2D0BWP U616 ( .A1(\ML_int[8][170] ), .A2(n22), .Z(\ML_int[10][170] ) );
  NR2D0BWP U617 ( .A1(n5), .A2(n164), .ZN(\ML_int[10][16] ) );
  CKND2D0BWP U618 ( .A1(\ML_int[6][16] ), .A2(n107), .ZN(n164) );
  INR2D0BWP U619 ( .A1(\ML_int[5][16] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][16] ) );
  AN2D0BWP U620 ( .A1(\ML_int[8][169] ), .A2(n22), .Z(\ML_int[10][169] ) );
  AN2D0BWP U621 ( .A1(\ML_int[8][168] ), .A2(n22), .Z(\ML_int[10][168] ) );
  AN2D0BWP U622 ( .A1(\ML_int[8][167] ), .A2(n22), .Z(\ML_int[10][167] ) );
  AN2D0BWP U623 ( .A1(\ML_int[8][166] ), .A2(n22), .Z(\ML_int[10][166] ) );
  AN2D0BWP U624 ( .A1(\ML_int[8][165] ), .A2(n22), .Z(\ML_int[10][165] ) );
  AN2D0BWP U625 ( .A1(\ML_int[8][164] ), .A2(n23), .Z(\ML_int[10][164] ) );
  AN2D0BWP U626 ( .A1(\ML_int[8][163] ), .A2(n23), .Z(\ML_int[10][163] ) );
  AN2D0BWP U627 ( .A1(\ML_int[8][162] ), .A2(n23), .Z(\ML_int[10][162] ) );
  AN2D0BWP U628 ( .A1(\ML_int[8][161] ), .A2(n23), .Z(\ML_int[10][161] ) );
  AN2D0BWP U629 ( .A1(\ML_int[8][160] ), .A2(n23), .Z(\ML_int[10][160] ) );
  NR2D0BWP U630 ( .A1(n5), .A2(n165), .ZN(\ML_int[10][15] ) );
  CKND2D0BWP U631 ( .A1(\ML_int[6][15] ), .A2(n107), .ZN(n165) );
  INR2D0BWP U632 ( .A1(\ML_int[5][15] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][15] ) );
  INR2D0BWP U633 ( .A1(A[15]), .B1(\temp_int_SH[4] ), .ZN(\ML_int[5][15] ) );
  AN2D0BWP U634 ( .A1(\ML_int[8][159] ), .A2(n23), .Z(\ML_int[10][159] ) );
  AN2D0BWP U635 ( .A1(\ML_int[8][158] ), .A2(n23), .Z(\ML_int[10][158] ) );
  AN2D0BWP U636 ( .A1(\ML_int[8][157] ), .A2(n23), .Z(\ML_int[10][157] ) );
  AN2D0BWP U637 ( .A1(\ML_int[8][156] ), .A2(n23), .Z(\ML_int[10][156] ) );
  AN2D0BWP U638 ( .A1(\ML_int[8][155] ), .A2(n23), .Z(\ML_int[10][155] ) );
  AN2D0BWP U639 ( .A1(\ML_int[8][154] ), .A2(n23), .Z(\ML_int[10][154] ) );
  AN2D0BWP U640 ( .A1(\ML_int[8][153] ), .A2(n23), .Z(\ML_int[10][153] ) );
  AN2D0BWP U641 ( .A1(\ML_int[8][152] ), .A2(n23), .Z(\ML_int[10][152] ) );
  AN2D0BWP U642 ( .A1(\ML_int[8][151] ), .A2(n24), .Z(\ML_int[10][151] ) );
  AN2D0BWP U643 ( .A1(\ML_int[8][150] ), .A2(n24), .Z(\ML_int[10][150] ) );
  NR2D0BWP U644 ( .A1(n5), .A2(n166), .ZN(\ML_int[10][14] ) );
  CKND2D0BWP U645 ( .A1(\ML_int[6][14] ), .A2(n107), .ZN(n166) );
  INR2D0BWP U646 ( .A1(\ML_int[5][14] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][14] ) );
  INR2D0BWP U647 ( .A1(A[14]), .B1(\temp_int_SH[4] ), .ZN(\ML_int[5][14] ) );
  AN2D0BWP U648 ( .A1(\ML_int[8][149] ), .A2(n24), .Z(\ML_int[10][149] ) );
  AN2D0BWP U649 ( .A1(\ML_int[8][148] ), .A2(n24), .Z(\ML_int[10][148] ) );
  AN2D0BWP U650 ( .A1(\ML_int[8][147] ), .A2(n24), .Z(\ML_int[10][147] ) );
  AN2D0BWP U651 ( .A1(\ML_int[8][146] ), .A2(n24), .Z(\ML_int[10][146] ) );
  AN2D0BWP U652 ( .A1(\ML_int[8][145] ), .A2(n24), .Z(\ML_int[10][145] ) );
  AN2D0BWP U653 ( .A1(\ML_int[8][144] ), .A2(n24), .Z(\ML_int[10][144] ) );
  AN2D0BWP U654 ( .A1(\ML_int[8][143] ), .A2(n24), .Z(\ML_int[10][143] ) );
  AN2D0BWP U655 ( .A1(\ML_int[8][142] ), .A2(n24), .Z(\ML_int[10][142] ) );
  AN2D0BWP U656 ( .A1(\ML_int[8][141] ), .A2(n24), .Z(\ML_int[10][141] ) );
  AN2D0BWP U657 ( .A1(\ML_int[8][140] ), .A2(n24), .Z(\ML_int[10][140] ) );
  NR2D0BWP U658 ( .A1(n6), .A2(n167), .ZN(\ML_int[10][13] ) );
  CKND2D0BWP U659 ( .A1(\ML_int[6][13] ), .A2(n107), .ZN(n167) );
  INR2D0BWP U660 ( .A1(\ML_int[5][13] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][13] ) );
  INR2D0BWP U661 ( .A1(A[13]), .B1(\temp_int_SH[4] ), .ZN(\ML_int[5][13] ) );
  AN2D0BWP U662 ( .A1(\ML_int[8][139] ), .A2(n24), .Z(\ML_int[10][139] ) );
  AN2D0BWP U663 ( .A1(\ML_int[8][138] ), .A2(n25), .Z(\ML_int[10][138] ) );
  AN2D0BWP U664 ( .A1(\ML_int[8][137] ), .A2(n25), .Z(\ML_int[10][137] ) );
  AN2D0BWP U665 ( .A1(\ML_int[8][136] ), .A2(n25), .Z(\ML_int[10][136] ) );
  AN2D0BWP U666 ( .A1(\ML_int[8][135] ), .A2(n25), .Z(\ML_int[10][135] ) );
  AN2D0BWP U667 ( .A1(\ML_int[8][134] ), .A2(n25), .Z(\ML_int[10][134] ) );
  AN2D0BWP U668 ( .A1(\ML_int[8][133] ), .A2(n25), .Z(\ML_int[10][133] ) );
  AN2D0BWP U669 ( .A1(\ML_int[8][132] ), .A2(n25), .Z(\ML_int[10][132] ) );
  AN2D0BWP U670 ( .A1(\ML_int[8][131] ), .A2(n25), .Z(\ML_int[10][131] ) );
  AN2D0BWP U671 ( .A1(\ML_int[8][130] ), .A2(n25), .Z(\ML_int[10][130] ) );
  NR2D0BWP U672 ( .A1(n6), .A2(n168), .ZN(\ML_int[10][12] ) );
  CKND2D0BWP U673 ( .A1(\ML_int[6][12] ), .A2(n107), .ZN(n168) );
  INR2D0BWP U674 ( .A1(\ML_int[5][12] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][12] ) );
  INR2D0BWP U675 ( .A1(A[12]), .B1(\temp_int_SH[4] ), .ZN(\ML_int[5][12] ) );
  AN2D0BWP U676 ( .A1(\ML_int[8][129] ), .A2(n25), .Z(\ML_int[10][129] ) );
  AN2D0BWP U677 ( .A1(\ML_int[8][128] ), .A2(n25), .Z(\ML_int[10][128] ) );
  INR2D0BWP U678 ( .A1(\ML_int[7][127] ), .B1(n6), .ZN(\ML_int[10][127] ) );
  INR2D0BWP U679 ( .A1(\ML_int[7][126] ), .B1(n6), .ZN(\ML_int[10][126] ) );
  INR2D0BWP U680 ( .A1(\ML_int[7][125] ), .B1(n6), .ZN(\ML_int[10][125] ) );
  INR2D0BWP U681 ( .A1(\ML_int[7][124] ), .B1(n6), .ZN(\ML_int[10][124] ) );
  INR2D0BWP U682 ( .A1(\ML_int[7][123] ), .B1(n6), .ZN(\ML_int[10][123] ) );
  INR2D0BWP U683 ( .A1(\ML_int[7][122] ), .B1(n6), .ZN(\ML_int[10][122] ) );
  INR2D0BWP U684 ( .A1(\ML_int[7][121] ), .B1(n6), .ZN(\ML_int[10][121] ) );
  INR2D0BWP U685 ( .A1(\ML_int[7][120] ), .B1(n6), .ZN(\ML_int[10][120] ) );
  NR2D0BWP U686 ( .A1(n6), .A2(n169), .ZN(\ML_int[10][11] ) );
  CKND2D0BWP U687 ( .A1(\ML_int[6][11] ), .A2(n107), .ZN(n169) );
  INR2D0BWP U688 ( .A1(\ML_int[5][11] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][11] ) );
  INR2D0BWP U689 ( .A1(A[11]), .B1(\temp_int_SH[4] ), .ZN(\ML_int[5][11] ) );
  INR2D0BWP U690 ( .A1(\ML_int[7][119] ), .B1(n6), .ZN(\ML_int[10][119] ) );
  INR2D0BWP U691 ( .A1(\ML_int[7][118] ), .B1(n7), .ZN(\ML_int[10][118] ) );
  INR2D0BWP U692 ( .A1(\ML_int[7][117] ), .B1(n7), .ZN(\ML_int[10][117] ) );
  INR2D0BWP U693 ( .A1(\ML_int[7][116] ), .B1(n7), .ZN(\ML_int[10][116] ) );
  INR2D0BWP U694 ( .A1(\ML_int[7][115] ), .B1(n7), .ZN(\ML_int[10][115] ) );
  INR2D0BWP U695 ( .A1(\ML_int[7][114] ), .B1(n7), .ZN(\ML_int[10][114] ) );
  INR2D0BWP U696 ( .A1(\ML_int[7][113] ), .B1(n7), .ZN(\ML_int[10][113] ) );
  INR2D0BWP U697 ( .A1(\ML_int[7][112] ), .B1(n7), .ZN(\ML_int[10][112] ) );
  INR2D0BWP U698 ( .A1(\ML_int[7][111] ), .B1(n7), .ZN(\ML_int[10][111] ) );
  INR2D0BWP U699 ( .A1(\ML_int[7][110] ), .B1(n7), .ZN(\ML_int[10][110] ) );
  NR2D0BWP U700 ( .A1(n6), .A2(n170), .ZN(\ML_int[10][10] ) );
  CKND2D0BWP U701 ( .A1(\ML_int[6][10] ), .A2(n107), .ZN(n170) );
  INR2D0BWP U702 ( .A1(\ML_int[5][10] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][10] ) );
  INR2D0BWP U703 ( .A1(A[10]), .B1(\temp_int_SH[4] ), .ZN(\ML_int[5][10] ) );
  INR2D0BWP U704 ( .A1(\ML_int[7][109] ), .B1(n7), .ZN(\ML_int[10][109] ) );
  INR2D0BWP U705 ( .A1(\ML_int[7][108] ), .B1(n7), .ZN(\ML_int[10][108] ) );
  INR2D0BWP U706 ( .A1(\ML_int[7][107] ), .B1(n7), .ZN(\ML_int[10][107] ) );
  INR2D0BWP U707 ( .A1(\ML_int[7][106] ), .B1(n7), .ZN(\ML_int[10][106] ) );
  INR2D0BWP U708 ( .A1(\ML_int[7][105] ), .B1(n8), .ZN(\ML_int[10][105] ) );
  INR2D0BWP U709 ( .A1(\ML_int[7][104] ), .B1(n8), .ZN(\ML_int[10][104] ) );
  INR2D0BWP U710 ( .A1(\ML_int[7][103] ), .B1(n8), .ZN(\ML_int[10][103] ) );
  INR2D0BWP U711 ( .A1(\ML_int[7][102] ), .B1(n9), .ZN(\ML_int[10][102] ) );
  INR2D0BWP U712 ( .A1(\ML_int[7][101] ), .B1(n10), .ZN(\ML_int[10][101] ) );
  INR2D0BWP U713 ( .A1(\ML_int[7][100] ), .B1(n11), .ZN(\ML_int[10][100] ) );
  NR2D0BWP U714 ( .A1(n4), .A2(n171), .ZN(\ML_int[10][0] ) );
  CKND2D0BWP U715 ( .A1(\ML_int[6][0] ), .A2(n107), .ZN(n171) );
  INR2D0BWP U716 ( .A1(\ML_int[5][0] ), .B1(\temp_int_SH[5] ), .ZN(
        \ML_int[6][0] ) );
  INR2D0BWP U717 ( .A1(\ML_int[4][0] ), .B1(\temp_int_SH[4] ), .ZN(
        \ML_int[5][0] ) );
  CKND2D0BWP U718 ( .A1(n25), .A2(n41), .ZN(n172) );
  NR2D0BWP U719 ( .A1(SH[9]), .A2(SH[8]), .ZN(n173) );
endmodule


module CVP14_DW01_inc_1 ( A, SUM );
  input [26:0] A;
  output [26:0] SUM;
  wire   n1, n2, n3, n4;
  wire   [26:2] carry;

  HA1D0BWP U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(SUM[26]), .S(SUM[25]) );
  HA1D0BWP U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  HA1D0BWP U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  HA1D0BWP U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  HA1D0BWP U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  HA1D0BWP U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  HA1D0BWP U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  HA1D0BWP U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  HA1D0BWP U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  HA1D0BWP U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  HA1D0BWP U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  HA1D0BWP U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  HA1D0BWP U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  NR4D0BWP U1 ( .A1(n1), .A2(n2), .A3(n3), .A4(n4), .ZN(carry[13]) );
  ND3D0BWP U2 ( .A1(A[8]), .A2(A[7]), .A3(A[9]), .ZN(n4) );
  ND3D0BWP U3 ( .A1(A[5]), .A2(A[4]), .A3(A[6]), .ZN(n3) );
  ND3D0BWP U4 ( .A1(A[2]), .A2(A[1]), .A3(A[3]), .ZN(n2) );
  ND4D0BWP U5 ( .A1(A[12]), .A2(A[11]), .A3(A[10]), .A4(A[0]), .ZN(n1) );
endmodule


module CVP14_DW01_ash_3 ( A, DATA_TC, SH, SH_TC, B );
  input [12:0] A;
  input [3:0] SH;
  output [12:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][12] , \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] ,
         \ML_int[1][8] , \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] ,
         \ML_int[1][4] , \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] ,
         \ML_int[1][0] , \ML_int[2][12] , \ML_int[2][11] , \ML_int[2][10] ,
         \ML_int[2][9] , \ML_int[2][8] , \ML_int[2][7] , \ML_int[2][6] ,
         \ML_int[2][5] , \ML_int[2][4] , \ML_int[2][3] , \ML_int[2][2] ,
         \ML_int[3][12] , \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] ,
         \ML_int[3][8] , \ML_int[3][5] , \ML_int[3][4] , \ML_int[3][3] ,
         \ML_int[3][2] , \ML_int[3][1] , \ML_int[3][0] , \ML_int[4][12] ,
         \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] ,
         \ML_int[4][7] , \ML_int[4][6] , \ML_int[4][5] , \ML_int[4][4] ,
         \ML_int[4][3] , \ML_int[4][2] , \ML_int[4][1] , \ML_int[4][0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10;
  assign B[12] = \ML_int[4][12] ;
  assign B[11] = \ML_int[4][11] ;
  assign B[10] = \ML_int[4][10] ;
  assign B[9] = \ML_int[4][9] ;
  assign B[8] = \ML_int[4][8] ;
  assign B[7] = \ML_int[4][7] ;
  assign B[6] = \ML_int[4][6] ;
  assign B[5] = \ML_int[4][5] ;
  assign B[4] = \ML_int[4][4] ;
  assign B[3] = \ML_int[4][3] ;
  assign B[2] = \ML_int[4][2] ;
  assign B[1] = \ML_int[4][1] ;
  assign B[0] = \ML_int[4][0] ;

  MUX2D0BWP M1_0_11 ( .I0(A[11]), .I1(A[10]), .S(SH[0]), .Z(\ML_int[1][11] )
         );
  MUX2D0BWP M1_1_11 ( .I0(\ML_int[1][11] ), .I1(\ML_int[1][9] ), .S(SH[1]), 
        .Z(\ML_int[2][11] ) );
  MUX2D0BWP M1_0_12 ( .I0(A[12]), .I1(A[11]), .S(SH[0]), .Z(\ML_int[1][12] )
         );
  MUX2D0BWP M1_0_10 ( .I0(A[10]), .I1(A[9]), .S(SH[0]), .Z(\ML_int[1][10] ) );
  MUX2D0BWP M1_0_8 ( .I0(A[8]), .I1(A[7]), .S(SH[0]), .Z(\ML_int[1][8] ) );
  MUX2D0BWP M1_0_6 ( .I0(A[6]), .I1(A[5]), .S(SH[0]), .Z(\ML_int[1][6] ) );
  MUX2D0BWP M1_0_9 ( .I0(A[9]), .I1(A[8]), .S(SH[0]), .Z(\ML_int[1][9] ) );
  MUX2D0BWP M1_0_7 ( .I0(A[7]), .I1(A[6]), .S(SH[0]), .Z(\ML_int[1][7] ) );
  MUX2D0BWP M1_0_5 ( .I0(A[5]), .I1(A[4]), .S(SH[0]), .Z(\ML_int[1][5] ) );
  MUX2D0BWP M1_0_4 ( .I0(A[4]), .I1(A[3]), .S(SH[0]), .Z(\ML_int[1][4] ) );
  MUX2D0BWP M1_0_3 ( .I0(A[3]), .I1(A[2]), .S(SH[0]), .Z(\ML_int[1][3] ) );
  MUX2D0BWP M1_0_2 ( .I0(A[2]), .I1(A[1]), .S(SH[0]), .Z(\ML_int[1][2] ) );
  MUX2D0BWP M1_1_12 ( .I0(\ML_int[1][12] ), .I1(\ML_int[1][10] ), .S(SH[1]), 
        .Z(\ML_int[2][12] ) );
  MUX2D0BWP M1_2_12 ( .I0(\ML_int[2][12] ), .I1(\ML_int[2][8] ), .S(SH[2]), 
        .Z(\ML_int[3][12] ) );
  MUX2D1BWP M1_3_12 ( .I0(\ML_int[3][12] ), .I1(\ML_int[3][4] ), .S(SH[3]), 
        .Z(\ML_int[4][12] ) );
  MUX2D0BWP M1_2_10 ( .I0(\ML_int[2][10] ), .I1(\ML_int[2][6] ), .S(SH[2]), 
        .Z(\ML_int[3][10] ) );
  MUX2D1BWP M1_3_10 ( .I0(\ML_int[3][10] ), .I1(\ML_int[3][2] ), .S(SH[3]), 
        .Z(\ML_int[4][10] ) );
  MUX2D0BWP M1_2_9 ( .I0(\ML_int[2][9] ), .I1(\ML_int[2][5] ), .S(SH[2]), .Z(
        \ML_int[3][9] ) );
  MUX2D1BWP M1_3_9 ( .I0(\ML_int[3][9] ), .I1(\ML_int[3][1] ), .S(SH[3]), .Z(
        \ML_int[4][9] ) );
  MUX2D0BWP M1_2_5 ( .I0(\ML_int[2][5] ), .I1(n5), .S(SH[2]), .Z(
        \ML_int[3][5] ) );
  MUX2D0BWP M1_2_11 ( .I0(\ML_int[2][11] ), .I1(\ML_int[2][7] ), .S(SH[2]), 
        .Z(\ML_int[3][11] ) );
  MUX2D1BWP M1_3_11 ( .I0(\ML_int[3][11] ), .I1(\ML_int[3][3] ), .S(SH[3]), 
        .Z(\ML_int[4][11] ) );
  MUX2D0BWP M1_2_8 ( .I0(\ML_int[2][8] ), .I1(\ML_int[2][4] ), .S(SH[2]), .Z(
        \ML_int[3][8] ) );
  MUX2D1BWP M1_3_8 ( .I0(\ML_int[3][8] ), .I1(\ML_int[3][0] ), .S(SH[3]), .Z(
        \ML_int[4][8] ) );
  MUX2D0BWP M1_1_10 ( .I0(\ML_int[1][10] ), .I1(\ML_int[1][8] ), .S(SH[1]), 
        .Z(\ML_int[2][10] ) );
  MUX2D0BWP M1_1_9 ( .I0(\ML_int[1][9] ), .I1(\ML_int[1][7] ), .S(SH[1]), .Z(
        \ML_int[2][9] ) );
  MUX2D0BWP M1_1_8 ( .I0(\ML_int[1][8] ), .I1(\ML_int[1][6] ), .S(SH[1]), .Z(
        \ML_int[2][8] ) );
  MUX2D0BWP M1_1_7 ( .I0(\ML_int[1][7] ), .I1(\ML_int[1][5] ), .S(SH[1]), .Z(
        \ML_int[2][7] ) );
  MUX2D0BWP M1_1_6 ( .I0(\ML_int[1][6] ), .I1(\ML_int[1][4] ), .S(SH[1]), .Z(
        \ML_int[2][6] ) );
  MUX2D0BWP M1_1_5 ( .I0(\ML_int[1][5] ), .I1(\ML_int[1][3] ), .S(SH[1]), .Z(
        \ML_int[2][5] ) );
  MUX2D0BWP M1_1_4 ( .I0(\ML_int[1][4] ), .I1(\ML_int[1][2] ), .S(SH[1]), .Z(
        \ML_int[2][4] ) );
  MUX2D0BWP M1_0_1 ( .I0(A[1]), .I1(A[0]), .S(SH[0]), .Z(\ML_int[1][1] ) );
  MUX2D0BWP M1_1_3 ( .I0(\ML_int[1][3] ), .I1(\ML_int[1][1] ), .S(SH[1]), .Z(
        \ML_int[2][3] ) );
  MUX2D0BWP M1_1_2 ( .I0(\ML_int[1][2] ), .I1(\ML_int[1][0] ), .S(SH[1]), .Z(
        \ML_int[2][2] ) );
  MUX2D0BWP M1_2_4 ( .I0(\ML_int[2][4] ), .I1(n3), .S(SH[2]), .Z(
        \ML_int[3][4] ) );
  OR2D0BWP U3 ( .A1(SH[3]), .A2(SH[2]), .Z(n8) );
  INVD1BWP U4 ( .I(SH[1]), .ZN(n7) );
  INVD1BWP U5 ( .I(\ML_int[2][2] ), .ZN(n4) );
  INVD1BWP U6 ( .I(\ML_int[2][3] ), .ZN(n6) );
  INVD1BWP U7 ( .I(n10), .ZN(n3) );
  NR2XD0BWP U8 ( .A1(n1), .A2(SH[3]), .ZN(\ML_int[4][6] ) );
  MUX2ND0BWP U9 ( .I0(\ML_int[2][6] ), .I1(\ML_int[2][2] ), .S(SH[2]), .ZN(n1)
         );
  NR2XD0BWP U10 ( .A1(n2), .A2(SH[3]), .ZN(\ML_int[4][7] ) );
  MUX2ND0BWP U11 ( .I0(\ML_int[2][7] ), .I1(\ML_int[2][3] ), .S(SH[2]), .ZN(n2) );
  INVD1BWP U12 ( .I(n9), .ZN(n5) );
  INR2D0BWP U13 ( .A1(\ML_int[3][5] ), .B1(SH[3]), .ZN(\ML_int[4][5] ) );
  INR2D0BWP U14 ( .A1(\ML_int[3][4] ), .B1(SH[3]), .ZN(\ML_int[4][4] ) );
  NR2D0BWP U15 ( .A1(n8), .A2(n6), .ZN(\ML_int[4][3] ) );
  NR2D0BWP U16 ( .A1(n8), .A2(n4), .ZN(\ML_int[4][2] ) );
  NR2D0BWP U17 ( .A1(n8), .A2(n9), .ZN(\ML_int[4][1] ) );
  NR2D0BWP U18 ( .A1(n8), .A2(n10), .ZN(\ML_int[4][0] ) );
  NR2D0BWP U19 ( .A1(SH[2]), .A2(n6), .ZN(\ML_int[3][3] ) );
  NR2D0BWP U20 ( .A1(SH[2]), .A2(n4), .ZN(\ML_int[3][2] ) );
  NR2D0BWP U21 ( .A1(SH[2]), .A2(n9), .ZN(\ML_int[3][1] ) );
  NR2D0BWP U22 ( .A1(SH[2]), .A2(n10), .ZN(\ML_int[3][0] ) );
  CKND2D0BWP U23 ( .A1(\ML_int[1][1] ), .A2(n7), .ZN(n9) );
  CKND2D0BWP U24 ( .A1(\ML_int[1][0] ), .A2(n7), .ZN(n10) );
  INR2D0BWP U25 ( .A1(A[0]), .B1(SH[0]), .ZN(\ML_int[1][0] ) );
endmodule


module CVP14_DW01_addsub_1 ( A, B, CI, ADD_SUB, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [16:0] carry;
  wire   [15:0] B_AS;
  assign carry[0] = ADD_SUB;

  FA1D0BWP U1_4 ( .A(A[4]), .B(B_AS[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FA1D0BWP U1_3 ( .A(A[3]), .B(B_AS[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FA1D0BWP U1_2 ( .A(A[2]), .B(B_AS[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FA1D0BWP U1_1 ( .A(A[1]), .B(B_AS[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  XOR3D0BWP U1_15 ( .A1(A[15]), .A2(carry[0]), .A3(carry[15]), .Z(SUM[15]) );
  FA1D0BWP U1_0 ( .A(A[0]), .B(B_AS[0]), .CI(carry[0]), .CO(carry[1]), .S(
        SUM[0]) );
  FA1D0BWP U1_14 ( .A(A[14]), .B(carry[0]), .CI(carry[14]), .CO(carry[15]), 
        .S(SUM[14]) );
  FA1D0BWP U1_13 ( .A(A[13]), .B(carry[0]), .CI(carry[13]), .CO(carry[14]), 
        .S(SUM[13]) );
  FA1D0BWP U1_12 ( .A(A[12]), .B(carry[0]), .CI(carry[12]), .CO(carry[13]), 
        .S(SUM[12]) );
  FA1D0BWP U1_11 ( .A(A[11]), .B(carry[0]), .CI(carry[11]), .CO(carry[12]), 
        .S(SUM[11]) );
  FA1D0BWP U1_10 ( .A(A[10]), .B(carry[0]), .CI(carry[10]), .CO(carry[11]), 
        .S(SUM[10]) );
  FA1D0BWP U1_9 ( .A(A[9]), .B(carry[0]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FA1D0BWP U1_8 ( .A(A[8]), .B(carry[0]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  FA1D0BWP U1_7 ( .A(A[7]), .B(carry[0]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  FA1D0BWP U1_6 ( .A(A[6]), .B(carry[0]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FA1D0BWP U1_5 ( .A(A[5]), .B(carry[0]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  CKXOR2D0BWP U1 ( .A1(B[4]), .A2(carry[0]), .Z(B_AS[4]) );
  CKXOR2D0BWP U2 ( .A1(B[3]), .A2(carry[0]), .Z(B_AS[3]) );
  CKXOR2D0BWP U3 ( .A1(B[2]), .A2(carry[0]), .Z(B_AS[2]) );
  CKXOR2D0BWP U4 ( .A1(B[1]), .A2(carry[0]), .Z(B_AS[1]) );
  CKXOR2D0BWP U5 ( .A1(B[0]), .A2(carry[0]), .Z(B_AS[0]) );
endmodule


module CVP14_DW01_addsub_2 ( A, B, CI, ADD_SUB, SUM, CO );
  input [26:0] A;
  input [26:0] B;
  output [26:0] SUM;
  input CI, ADD_SUB;
  output CO;
  wire   n1, n2;
  wire   [27:0] carry;
  wire   [26:0] B_AS;
  assign carry[0] = ADD_SUB;

  FA1D0BWP U1_16 ( .A(A[16]), .B(B_AS[16]), .CI(carry[16]), .CO(carry[17]), 
        .S(SUM[16]) );
  FA1D0BWP U1_17 ( .A(A[17]), .B(B_AS[17]), .CI(carry[17]), .CO(carry[18]), 
        .S(SUM[17]) );
  FA1D0BWP U1_21 ( .A(A[21]), .B(B_AS[21]), .CI(carry[21]), .CO(carry[22]), 
        .S(SUM[21]) );
  FA1D0BWP U1_19 ( .A(A[19]), .B(B_AS[19]), .CI(carry[19]), .CO(carry[20]), 
        .S(SUM[19]) );
  FA1D0BWP U1_15 ( .A(A[15]), .B(B_AS[15]), .CI(carry[15]), .CO(carry[16]), 
        .S(SUM[15]) );
  FA1D0BWP U1_24 ( .A(A[24]), .B(B_AS[24]), .CI(carry[24]), .CO(carry[25]), 
        .S(SUM[24]) );
  FA1D0BWP U1_20 ( .A(A[20]), .B(B_AS[20]), .CI(carry[20]), .CO(carry[21]), 
        .S(SUM[20]) );
  FA1D0BWP U1_18 ( .A(A[18]), .B(B_AS[18]), .CI(carry[18]), .CO(carry[19]), 
        .S(SUM[18]) );
  FA1D0BWP U1_23 ( .A(A[23]), .B(B_AS[23]), .CI(carry[23]), .CO(carry[24]), 
        .S(SUM[23]) );
  FA1D0BWP U1_22 ( .A(A[22]), .B(B_AS[22]), .CI(carry[22]), .CO(carry[23]), 
        .S(SUM[22]) );
  FA1D0BWP U1_25 ( .A(A[25]), .B(B_AS[25]), .CI(carry[25]), .CO(carry[26]), 
        .S(SUM[25]) );
  INVD1BWP U1 ( .I(carry[14]), .ZN(n2) );
  INVD1BWP U2 ( .I(B_AS[14]), .ZN(n1) );
  XOR2D1BWP U3 ( .A1(carry[14]), .A2(B_AS[14]), .Z(SUM[14]) );
  AN2XD1BWP U4 ( .A1(B_AS[1]), .A2(carry[1]), .Z(carry[2]) );
  AN2XD1BWP U5 ( .A1(B_AS[2]), .A2(carry[2]), .Z(carry[3]) );
  AN2XD1BWP U6 ( .A1(B_AS[3]), .A2(carry[3]), .Z(carry[4]) );
  AN2XD1BWP U7 ( .A1(B_AS[4]), .A2(carry[4]), .Z(carry[5]) );
  AN2XD1BWP U8 ( .A1(B_AS[5]), .A2(carry[5]), .Z(carry[6]) );
  AN2XD1BWP U9 ( .A1(B_AS[6]), .A2(carry[6]), .Z(carry[7]) );
  AN2XD1BWP U10 ( .A1(B_AS[7]), .A2(carry[7]), .Z(carry[8]) );
  AN2XD1BWP U11 ( .A1(B_AS[8]), .A2(carry[8]), .Z(carry[9]) );
  AN2XD1BWP U12 ( .A1(B_AS[9]), .A2(carry[9]), .Z(carry[10]) );
  AN2XD1BWP U13 ( .A1(B_AS[10]), .A2(carry[10]), .Z(carry[11]) );
  AN2XD1BWP U14 ( .A1(B_AS[11]), .A2(carry[11]), .Z(carry[12]) );
  AN2XD1BWP U15 ( .A1(B_AS[12]), .A2(carry[12]), .Z(carry[13]) );
  AN2XD1BWP U16 ( .A1(B_AS[13]), .A2(carry[13]), .Z(carry[14]) );
  XOR2D1BWP U17 ( .A1(carry[13]), .A2(B_AS[13]), .Z(SUM[13]) );
  XOR2D1BWP U18 ( .A1(carry[5]), .A2(B_AS[5]), .Z(SUM[5]) );
  XOR2D1BWP U19 ( .A1(carry[9]), .A2(B_AS[9]), .Z(SUM[9]) );
  XOR2D1BWP U20 ( .A1(carry[1]), .A2(B_AS[1]), .Z(SUM[1]) );
  XOR2D1BWP U21 ( .A1(carry[6]), .A2(B_AS[6]), .Z(SUM[6]) );
  XOR2D1BWP U22 ( .A1(carry[10]), .A2(B_AS[10]), .Z(SUM[10]) );
  XOR2D1BWP U23 ( .A1(carry[2]), .A2(B_AS[2]), .Z(SUM[2]) );
  XOR2D1BWP U24 ( .A1(carry[7]), .A2(B_AS[7]), .Z(SUM[7]) );
  XOR2D1BWP U25 ( .A1(carry[11]), .A2(B_AS[11]), .Z(SUM[11]) );
  XOR2D1BWP U26 ( .A1(carry[3]), .A2(B_AS[3]), .Z(SUM[3]) );
  XOR2D1BWP U27 ( .A1(carry[8]), .A2(B_AS[8]), .Z(SUM[8]) );
  XOR2D1BWP U28 ( .A1(carry[12]), .A2(B_AS[12]), .Z(SUM[12]) );
  XOR2D1BWP U29 ( .A1(carry[4]), .A2(B_AS[4]), .Z(SUM[4]) );
  XOR2D1BWP U30 ( .A1(carry[0]), .A2(carry[26]), .Z(SUM[26]) );
  AN2XD1BWP U31 ( .A1(B_AS[0]), .A2(carry[0]), .Z(carry[1]) );
  CKXOR2D0BWP U32 ( .A1(carry[0]), .A2(B_AS[0]), .Z(SUM[0]) );
  NR2XD0BWP U33 ( .A1(n1), .A2(n2), .ZN(carry[15]) );
  CKXOR2D0BWP U34 ( .A1(B[9]), .A2(carry[0]), .Z(B_AS[9]) );
  CKXOR2D0BWP U35 ( .A1(B[8]), .A2(carry[0]), .Z(B_AS[8]) );
  CKXOR2D0BWP U36 ( .A1(B[7]), .A2(carry[0]), .Z(B_AS[7]) );
  CKXOR2D0BWP U37 ( .A1(B[6]), .A2(carry[0]), .Z(B_AS[6]) );
  CKXOR2D0BWP U38 ( .A1(B[5]), .A2(carry[0]), .Z(B_AS[5]) );
  CKXOR2D0BWP U39 ( .A1(B[4]), .A2(carry[0]), .Z(B_AS[4]) );
  CKXOR2D0BWP U40 ( .A1(B[3]), .A2(carry[0]), .Z(B_AS[3]) );
  CKXOR2D0BWP U41 ( .A1(B[2]), .A2(carry[0]), .Z(B_AS[2]) );
  CKXOR2D0BWP U42 ( .A1(B[25]), .A2(carry[0]), .Z(B_AS[25]) );
  CKXOR2D0BWP U43 ( .A1(B[24]), .A2(carry[0]), .Z(B_AS[24]) );
  CKXOR2D0BWP U44 ( .A1(B[23]), .A2(carry[0]), .Z(B_AS[23]) );
  CKXOR2D0BWP U45 ( .A1(B[22]), .A2(carry[0]), .Z(B_AS[22]) );
  CKXOR2D0BWP U46 ( .A1(B[21]), .A2(carry[0]), .Z(B_AS[21]) );
  CKXOR2D0BWP U47 ( .A1(B[20]), .A2(carry[0]), .Z(B_AS[20]) );
  CKXOR2D0BWP U48 ( .A1(B[1]), .A2(carry[0]), .Z(B_AS[1]) );
  CKXOR2D0BWP U49 ( .A1(B[19]), .A2(carry[0]), .Z(B_AS[19]) );
  CKXOR2D0BWP U50 ( .A1(B[18]), .A2(carry[0]), .Z(B_AS[18]) );
  CKXOR2D0BWP U51 ( .A1(B[17]), .A2(carry[0]), .Z(B_AS[17]) );
  CKXOR2D0BWP U52 ( .A1(B[16]), .A2(carry[0]), .Z(B_AS[16]) );
  CKXOR2D0BWP U53 ( .A1(B[15]), .A2(carry[0]), .Z(B_AS[15]) );
  CKXOR2D0BWP U54 ( .A1(B[14]), .A2(carry[0]), .Z(B_AS[14]) );
  CKXOR2D0BWP U55 ( .A1(B[13]), .A2(carry[0]), .Z(B_AS[13]) );
  CKXOR2D0BWP U56 ( .A1(B[12]), .A2(carry[0]), .Z(B_AS[12]) );
  CKXOR2D0BWP U57 ( .A1(B[11]), .A2(carry[0]), .Z(B_AS[11]) );
  CKXOR2D0BWP U58 ( .A1(B[10]), .A2(carry[0]), .Z(B_AS[10]) );
  CKXOR2D0BWP U59 ( .A1(B[0]), .A2(carry[0]), .Z(B_AS[0]) );
endmodule


module CVP14_DW_rash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [25:0] A;
  input [4:0] SH;
  output [25:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76;

  INVD1BWP U3 ( .I(n65), .ZN(n26) );
  INVD1BWP U4 ( .I(n66), .ZN(n25) );
  INVD1BWP U5 ( .I(n41), .ZN(n15) );
  INVD1BWP U6 ( .I(n37), .ZN(n2) );
  INVD1BWP U7 ( .I(n36), .ZN(n17) );
  INVD1BWP U8 ( .I(n40), .ZN(n1) );
  INVD1BWP U9 ( .I(n34), .ZN(n20) );
  INVD1BWP U10 ( .I(SH[0]), .ZN(n28) );
  INVD1BWP U11 ( .I(A[25]), .ZN(n29) );
  INVD1BWP U12 ( .I(n56), .ZN(n10) );
  INVD1BWP U13 ( .I(n38), .ZN(n11) );
  INVD1BWP U14 ( .I(n69), .ZN(n5) );
  INVD1BWP U15 ( .I(n57), .ZN(n23) );
  INVD1BWP U16 ( .I(n58), .ZN(n22) );
  INVD1BWP U17 ( .I(n67), .ZN(n18) );
  INVD1BWP U18 ( .I(SH[1]), .ZN(n27) );
  INVD1BWP U19 ( .I(n52), .ZN(n19) );
  INVD1BWP U20 ( .I(SH[4]), .ZN(n21) );
  INVD1BWP U21 ( .I(SH[2]), .ZN(n24) );
  INVD1BWP U22 ( .I(A[21]), .ZN(n12) );
  INVD1BWP U23 ( .I(A[24]), .ZN(n16) );
  INVD1BWP U24 ( .I(A[23]), .ZN(n14) );
  INVD1BWP U25 ( .I(A[22]), .ZN(n13) );
  INVD1BWP U26 ( .I(A[17]), .ZN(n6) );
  INVD1BWP U27 ( .I(A[16]), .ZN(n4) );
  INVD1BWP U28 ( .I(A[20]), .ZN(n9) );
  INVD1BWP U29 ( .I(A[19]), .ZN(n8) );
  INVD1BWP U30 ( .I(A[18]), .ZN(n7) );
  INVD1BWP U31 ( .I(A[15]), .ZN(n3) );
  OAI221D0BWP U32 ( .A1(n30), .A2(n31), .B1(n11), .B2(n32), .C(n33), .ZN(B[9])
         );
  AOI22D0BWP U33 ( .A1(n34), .A2(n35), .B1(n36), .B2(n37), .ZN(n33) );
  OAI221D0BWP U34 ( .A1(n5), .A2(n31), .B1(n10), .B2(n32), .C(n39), .ZN(B[8])
         );
  AOI22D0BWP U35 ( .A1(n40), .A2(n36), .B1(n34), .B2(n41), .ZN(n39) );
  OAI222D0BWP U36 ( .A1(n42), .A2(n31), .B1(n43), .B2(n20), .C1(n44), .C2(n32), 
        .ZN(B[7]) );
  OAI222D0BWP U37 ( .A1(n45), .A2(n31), .B1(n46), .B2(n20), .C1(n47), .C2(n32), 
        .ZN(B[6]) );
  NR2D0BWP U38 ( .A1(n21), .A2(n23), .ZN(n34) );
  OAI21D0BWP U39 ( .A1(n30), .A2(n32), .B(n48), .ZN(B[5]) );
  OA32D0BWP U40 ( .A1(n49), .A2(SH[3]), .A3(n21), .B1(n31), .B2(n2), .Z(n48)
         );
  OAI22D0BWP U41 ( .A1(n50), .A2(n21), .B1(n51), .B2(n52), .ZN(B[4]) );
  OAI22D0BWP U42 ( .A1(n53), .A2(n21), .B1(n42), .B2(n32), .ZN(B[3]) );
  OAI22D0BWP U43 ( .A1(n54), .A2(n21), .B1(n45), .B2(n32), .ZN(B[2]) );
  INR2D0BWP U44 ( .A1(n35), .B1(n55), .ZN(B[25]) );
  NR2D0BWP U45 ( .A1(n15), .A2(n55), .ZN(B[24]) );
  NR2D0BWP U46 ( .A1(n43), .A2(n55), .ZN(B[23]) );
  NR2D0BWP U47 ( .A1(n46), .A2(n55), .ZN(B[22]) );
  NR2D0BWP U48 ( .A1(n49), .A2(n18), .ZN(B[21]) );
  NR2D0BWP U49 ( .A1(SH[4]), .A2(n50), .ZN(B[20]) );
  AOI22D0BWP U50 ( .A1(n56), .A2(n57), .B1(n41), .B2(n58), .ZN(n50) );
  OAI22D0BWP U51 ( .A1(n59), .A2(n21), .B1(n2), .B2(n32), .ZN(B[1]) );
  NR2D0BWP U52 ( .A1(SH[4]), .A2(n53), .ZN(B[19]) );
  OA22D1BWP U53 ( .A1(n44), .A2(n23), .B1(n43), .B2(n22), .Z(n53) );
  NR2D0BWP U54 ( .A1(SH[4]), .A2(n54), .ZN(B[18]) );
  OA22D1BWP U55 ( .A1(n47), .A2(n23), .B1(n46), .B2(n22), .Z(n54) );
  NR2D0BWP U56 ( .A1(SH[4]), .A2(n59), .ZN(B[17]) );
  OA21D0BWP U57 ( .A1(n30), .A2(n23), .B(n60), .Z(n59) );
  AOI32D0BWP U58 ( .A1(n35), .A2(n24), .A3(SH[3]), .B1(n58), .B2(n38), .ZN(n60) );
  NR2D0BWP U59 ( .A1(SH[4]), .A2(n61), .ZN(B[16]) );
  OAI222D0BWP U60 ( .A1(n44), .A2(n17), .B1(n42), .B2(n55), .C1(n43), .C2(n31), 
        .ZN(B[15]) );
  OAI222D0BWP U61 ( .A1(n47), .A2(n17), .B1(n45), .B2(n55), .C1(n46), .C2(n31), 
        .ZN(B[14]) );
  OAI222D0BWP U62 ( .A1(n30), .A2(n17), .B1(n2), .B2(n55), .C1(n49), .C2(n52), 
        .ZN(B[13]) );
  MUX2ND0BWP U63 ( .I0(n35), .I1(n38), .S(n24), .ZN(n49) );
  OAI221D0BWP U64 ( .A1(n62), .A2(n13), .B1(n63), .B2(n14), .C(n64), .ZN(n38)
         );
  AOI22D0BWP U65 ( .A1(A[24]), .A2(n65), .B1(A[21]), .B2(n66), .ZN(n64) );
  NR2D0BWP U66 ( .A1(n29), .A2(n25), .ZN(n35) );
  CKND2D0BWP U67 ( .A1(n67), .A2(n24), .ZN(n55) );
  OAI22D0BWP U68 ( .A1(n26), .A2(n4), .B1(n63), .B2(n3), .ZN(n37) );
  OA221D0BWP U69 ( .A1(n62), .A2(n7), .B1(n63), .B2(n8), .C(n68), .Z(n30) );
  AOI22D0BWP U70 ( .A1(A[20]), .A2(n65), .B1(A[17]), .B2(n66), .ZN(n68) );
  OAI222D0BWP U71 ( .A1(n15), .A2(n32), .B1(n10), .B2(n31), .C1(n51), .C2(n18), 
        .ZN(B[12]) );
  MUX2ND0BWP U72 ( .I0(n69), .I1(n40), .S(n24), .ZN(n51) );
  OAI222D0BWP U73 ( .A1(n44), .A2(n31), .B1(n42), .B2(n17), .C1(n43), .C2(n32), 
        .ZN(B[11]) );
  OA222D0BWP U74 ( .A1(n29), .A2(n63), .B1(n62), .B2(n16), .C1(n25), .C2(n14), 
        .Z(n43) );
  OA221D0BWP U75 ( .A1(n4), .A2(n62), .B1(n63), .B2(n6), .C(n70), .Z(n42) );
  AOI22D0BWP U76 ( .A1(A[18]), .A2(n65), .B1(A[15]), .B2(n66), .ZN(n70) );
  OA221D0BWP U77 ( .A1(n62), .A2(n9), .B1(n63), .B2(n12), .C(n71), .Z(n44) );
  AOI22D0BWP U78 ( .A1(A[22]), .A2(n65), .B1(A[19]), .B2(n66), .ZN(n71) );
  OAI222D0BWP U79 ( .A1(n47), .A2(n31), .B1(n45), .B2(n17), .C1(n46), .C2(n32), 
        .ZN(B[10]) );
  OA221D0BWP U80 ( .A1(n62), .A2(n14), .B1(n63), .B2(n16), .C(n72), .Z(n46) );
  AOI22D0BWP U81 ( .A1(n65), .A2(A[25]), .B1(A[22]), .B2(n66), .ZN(n72) );
  NR2D0BWP U82 ( .A1(n24), .A2(n18), .ZN(n36) );
  NR2D0BWP U83 ( .A1(SH[3]), .A2(SH[4]), .ZN(n67) );
  OA222D0BWP U84 ( .A1(n63), .A2(n4), .B1(n3), .B2(n62), .C1(n26), .C2(n6), 
        .Z(n45) );
  CKND2D0BWP U85 ( .A1(n19), .A2(n24), .ZN(n31) );
  OA221D0BWP U86 ( .A1(n62), .A2(n8), .B1(n63), .B2(n9), .C(n73), .Z(n47) );
  AOI22D0BWP U87 ( .A1(A[21]), .A2(n65), .B1(A[18]), .B2(n66), .ZN(n73) );
  OAI22D0BWP U88 ( .A1(n61), .A2(n21), .B1(n32), .B2(n1), .ZN(B[0]) );
  NR2D0BWP U89 ( .A1(n26), .A2(n3), .ZN(n40) );
  CKND2D0BWP U90 ( .A1(n19), .A2(SH[2]), .ZN(n32) );
  CKND2D0BWP U91 ( .A1(SH[3]), .A2(n21), .ZN(n52) );
  OA21D0BWP U92 ( .A1(n5), .A2(n23), .B(n74), .Z(n61) );
  AOI32D0BWP U93 ( .A1(n41), .A2(n24), .A3(SH[3]), .B1(n58), .B2(n56), .ZN(n74) );
  OAI221D0BWP U94 ( .A1(n62), .A2(n12), .B1(n63), .B2(n13), .C(n75), .ZN(n56)
         );
  AOI22D0BWP U95 ( .A1(A[23]), .A2(n65), .B1(A[20]), .B2(n66), .ZN(n75) );
  NR2D0BWP U96 ( .A1(n24), .A2(SH[3]), .ZN(n58) );
  OAI22D0BWP U97 ( .A1(n25), .A2(n16), .B1(n29), .B2(n62), .ZN(n41) );
  NR2D0BWP U98 ( .A1(SH[2]), .A2(SH[3]), .ZN(n57) );
  OAI221D0BWP U99 ( .A1(n62), .A2(n6), .B1(n63), .B2(n7), .C(n76), .ZN(n69) );
  AOI22D0BWP U100 ( .A1(A[19]), .A2(n65), .B1(A[16]), .B2(n66), .ZN(n76) );
  NR2D0BWP U101 ( .A1(SH[0]), .A2(SH[1]), .ZN(n66) );
  NR2D0BWP U102 ( .A1(n28), .A2(n27), .ZN(n65) );
  CKND2D0BWP U103 ( .A1(SH[1]), .A2(n28), .ZN(n63) );
  CKND2D0BWP U104 ( .A1(SH[0]), .A2(n27), .ZN(n62) );
endmodule


module CVP14_DW_rash_1 ( A, DATA_TC, SH, SH_TC, B );
  input [25:0] A;
  input [4:0] SH;
  output [25:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76;

  INVD1BWP U3 ( .I(n65), .ZN(n16) );
  INVD1BWP U4 ( .I(n66), .ZN(n11) );
  INVD1BWP U5 ( .I(n36), .ZN(n1) );
  INVD1BWP U6 ( .I(n34), .ZN(n4) );
  CKND0BWP U7 ( .I(SH[0]), .ZN(n18) );
  INVD1BWP U8 ( .I(n41), .ZN(n10) );
  INVD1BWP U9 ( .I(n37), .ZN(n14) );
  INVD1BWP U10 ( .I(n57), .ZN(n7) );
  INVD1BWP U11 ( .I(n58), .ZN(n6) );
  INVD1BWP U12 ( .I(n67), .ZN(n2) );
  INVD1BWP U13 ( .I(n40), .ZN(n15) );
  INVD1BWP U14 ( .I(SH[1]), .ZN(n17) );
  INVD1BWP U15 ( .I(n52), .ZN(n3) );
  INVD1BWP U16 ( .I(A[25]), .ZN(n20) );
  CKND0BWP U17 ( .I(SH[4]), .ZN(n5) );
  INVD1BWP U18 ( .I(n56), .ZN(n12) );
  INVD1BWP U19 ( .I(n38), .ZN(n13) );
  CKND0BWP U20 ( .I(SH[2]), .ZN(n8) );
  INVD1BWP U21 ( .I(n69), .ZN(n9) );
  INVD1BWP U22 ( .I(A[17]), .ZN(n28) );
  INVD1BWP U23 ( .I(A[15]), .ZN(n19) );
  INVD1BWP U24 ( .I(A[16]), .ZN(n29) );
  INVD1BWP U25 ( .I(A[24]), .ZN(n21) );
  INVD1BWP U26 ( .I(A[23]), .ZN(n22) );
  INVD1BWP U27 ( .I(A[21]), .ZN(n24) );
  INVD1BWP U28 ( .I(A[22]), .ZN(n23) );
  INVD1BWP U29 ( .I(A[20]), .ZN(n25) );
  INVD1BWP U30 ( .I(A[19]), .ZN(n26) );
  INVD1BWP U31 ( .I(A[18]), .ZN(n27) );
  OAI221D0BWP U32 ( .A1(n30), .A2(n31), .B1(n13), .B2(n32), .C(n33), .ZN(B[9])
         );
  AOI22D0BWP U33 ( .A1(n34), .A2(n35), .B1(n36), .B2(n37), .ZN(n33) );
  OAI221D0BWP U34 ( .A1(n9), .A2(n31), .B1(n12), .B2(n32), .C(n39), .ZN(B[8])
         );
  AOI22D0BWP U35 ( .A1(n40), .A2(n36), .B1(n34), .B2(n41), .ZN(n39) );
  OAI222D0BWP U36 ( .A1(n42), .A2(n31), .B1(n43), .B2(n4), .C1(n44), .C2(n32), 
        .ZN(B[7]) );
  OAI222D0BWP U37 ( .A1(n45), .A2(n31), .B1(n46), .B2(n4), .C1(n47), .C2(n32), 
        .ZN(B[6]) );
  NR2D0BWP U38 ( .A1(n5), .A2(n7), .ZN(n34) );
  OAI21D0BWP U39 ( .A1(n30), .A2(n32), .B(n48), .ZN(B[5]) );
  OA32D0BWP U40 ( .A1(n49), .A2(SH[3]), .A3(n5), .B1(n31), .B2(n14), .Z(n48)
         );
  OAI22D0BWP U41 ( .A1(n50), .A2(n5), .B1(n51), .B2(n52), .ZN(B[4]) );
  OAI22D0BWP U42 ( .A1(n53), .A2(n5), .B1(n42), .B2(n32), .ZN(B[3]) );
  OAI22D0BWP U43 ( .A1(n54), .A2(n5), .B1(n45), .B2(n32), .ZN(B[2]) );
  INR2D0BWP U44 ( .A1(n35), .B1(n55), .ZN(B[25]) );
  NR2D0BWP U45 ( .A1(n10), .A2(n55), .ZN(B[24]) );
  NR2D0BWP U46 ( .A1(n43), .A2(n55), .ZN(B[23]) );
  NR2D0BWP U47 ( .A1(n46), .A2(n55), .ZN(B[22]) );
  NR2D0BWP U48 ( .A1(n49), .A2(n2), .ZN(B[21]) );
  NR2D0BWP U49 ( .A1(SH[4]), .A2(n50), .ZN(B[20]) );
  AOI22D0BWP U50 ( .A1(n56), .A2(n57), .B1(n41), .B2(n58), .ZN(n50) );
  OAI22D0BWP U51 ( .A1(n59), .A2(n5), .B1(n14), .B2(n32), .ZN(B[1]) );
  NR2D0BWP U52 ( .A1(SH[4]), .A2(n53), .ZN(B[19]) );
  OA22D1BWP U53 ( .A1(n44), .A2(n7), .B1(n43), .B2(n6), .Z(n53) );
  NR2D0BWP U54 ( .A1(SH[4]), .A2(n54), .ZN(B[18]) );
  OA22D1BWP U55 ( .A1(n47), .A2(n7), .B1(n46), .B2(n6), .Z(n54) );
  NR2D0BWP U56 ( .A1(SH[4]), .A2(n59), .ZN(B[17]) );
  OA21D0BWP U57 ( .A1(n30), .A2(n7), .B(n60), .Z(n59) );
  AOI32D0BWP U58 ( .A1(n35), .A2(n8), .A3(SH[3]), .B1(n58), .B2(n38), .ZN(n60)
         );
  NR2D0BWP U59 ( .A1(SH[4]), .A2(n61), .ZN(B[16]) );
  OAI222D0BWP U60 ( .A1(n44), .A2(n1), .B1(n42), .B2(n55), .C1(n43), .C2(n31), 
        .ZN(B[15]) );
  OAI222D0BWP U61 ( .A1(n47), .A2(n1), .B1(n45), .B2(n55), .C1(n46), .C2(n31), 
        .ZN(B[14]) );
  OAI222D0BWP U62 ( .A1(n30), .A2(n1), .B1(n14), .B2(n55), .C1(n49), .C2(n52), 
        .ZN(B[13]) );
  MUX2ND0BWP U63 ( .I0(n35), .I1(n38), .S(n8), .ZN(n49) );
  OAI221D0BWP U64 ( .A1(n62), .A2(n23), .B1(n63), .B2(n22), .C(n64), .ZN(n38)
         );
  AOI22D0BWP U65 ( .A1(A[24]), .A2(n65), .B1(A[21]), .B2(n66), .ZN(n64) );
  NR2D0BWP U66 ( .A1(n20), .A2(n11), .ZN(n35) );
  CKND2D0BWP U67 ( .A1(n67), .A2(n8), .ZN(n55) );
  OAI22D0BWP U68 ( .A1(n16), .A2(n29), .B1(n63), .B2(n19), .ZN(n37) );
  OA221D0BWP U69 ( .A1(n62), .A2(n27), .B1(n63), .B2(n26), .C(n68), .Z(n30) );
  AOI22D0BWP U70 ( .A1(A[20]), .A2(n65), .B1(A[17]), .B2(n66), .ZN(n68) );
  OAI222D0BWP U71 ( .A1(n10), .A2(n32), .B1(n12), .B2(n31), .C1(n51), .C2(n2), 
        .ZN(B[12]) );
  MUX2ND0BWP U72 ( .I0(n69), .I1(n40), .S(n8), .ZN(n51) );
  OAI222D0BWP U73 ( .A1(n44), .A2(n31), .B1(n42), .B2(n1), .C1(n43), .C2(n32), 
        .ZN(B[11]) );
  OA222D0BWP U74 ( .A1(n20), .A2(n63), .B1(n62), .B2(n21), .C1(n11), .C2(n22), 
        .Z(n43) );
  OA221D0BWP U75 ( .A1(n29), .A2(n62), .B1(n63), .B2(n28), .C(n70), .Z(n42) );
  AOI22D0BWP U76 ( .A1(A[18]), .A2(n65), .B1(A[15]), .B2(n66), .ZN(n70) );
  OA221D0BWP U77 ( .A1(n62), .A2(n25), .B1(n63), .B2(n24), .C(n71), .Z(n44) );
  AOI22D0BWP U78 ( .A1(A[22]), .A2(n65), .B1(A[19]), .B2(n66), .ZN(n71) );
  OAI222D0BWP U79 ( .A1(n47), .A2(n31), .B1(n45), .B2(n1), .C1(n46), .C2(n32), 
        .ZN(B[10]) );
  OA221D0BWP U80 ( .A1(n62), .A2(n22), .B1(n63), .B2(n21), .C(n72), .Z(n46) );
  AOI22D0BWP U81 ( .A1(n65), .A2(A[25]), .B1(A[22]), .B2(n66), .ZN(n72) );
  NR2D0BWP U82 ( .A1(n8), .A2(n2), .ZN(n36) );
  NR2D0BWP U83 ( .A1(SH[3]), .A2(SH[4]), .ZN(n67) );
  OA222D0BWP U84 ( .A1(n63), .A2(n29), .B1(n19), .B2(n62), .C1(n16), .C2(n28), 
        .Z(n45) );
  CKND2D0BWP U85 ( .A1(n3), .A2(n8), .ZN(n31) );
  OA221D0BWP U86 ( .A1(n62), .A2(n26), .B1(n63), .B2(n25), .C(n73), .Z(n47) );
  AOI22D0BWP U87 ( .A1(A[21]), .A2(n65), .B1(A[18]), .B2(n66), .ZN(n73) );
  OAI22D0BWP U88 ( .A1(n61), .A2(n5), .B1(n32), .B2(n15), .ZN(B[0]) );
  NR2D0BWP U89 ( .A1(n16), .A2(n19), .ZN(n40) );
  CKND2D0BWP U90 ( .A1(n3), .A2(SH[2]), .ZN(n32) );
  CKND2D0BWP U91 ( .A1(SH[3]), .A2(n5), .ZN(n52) );
  OA21D0BWP U92 ( .A1(n9), .A2(n7), .B(n74), .Z(n61) );
  AOI32D0BWP U93 ( .A1(n41), .A2(n8), .A3(SH[3]), .B1(n58), .B2(n56), .ZN(n74)
         );
  OAI221D0BWP U94 ( .A1(n62), .A2(n24), .B1(n63), .B2(n23), .C(n75), .ZN(n56)
         );
  AOI22D0BWP U95 ( .A1(A[23]), .A2(n65), .B1(A[20]), .B2(n66), .ZN(n75) );
  NR2D0BWP U96 ( .A1(n8), .A2(SH[3]), .ZN(n58) );
  OAI22D0BWP U97 ( .A1(n11), .A2(n21), .B1(n20), .B2(n62), .ZN(n41) );
  NR2D0BWP U98 ( .A1(SH[2]), .A2(SH[3]), .ZN(n57) );
  OAI221D0BWP U99 ( .A1(n62), .A2(n28), .B1(n63), .B2(n27), .C(n76), .ZN(n69)
         );
  AOI22D0BWP U100 ( .A1(A[19]), .A2(n65), .B1(A[16]), .B2(n66), .ZN(n76) );
  NR2D0BWP U101 ( .A1(SH[0]), .A2(SH[1]), .ZN(n66) );
  NR2D0BWP U102 ( .A1(n18), .A2(n17), .ZN(n65) );
  CKND2D0BWP U103 ( .A1(SH[1]), .A2(n18), .ZN(n63) );
  CKND2D0BWP U104 ( .A1(SH[0]), .A2(n17), .ZN(n62) );
endmodule


module CVP14_DW01_ash_4 ( A, DATA_TC, SH, SH_TC, B );
  input [11:0] A;
  input [3:0] SH;
  output [11:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[3][11] , \ML_int[3][10] ,
         \ML_int[3][9] , \ML_int[3][8] , \ML_int[3][1] , \ML_int[3][0] ,
         \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] ,
         \ML_int[4][7] , \ML_int[4][6] , \ML_int[4][5] , \ML_int[4][4] ,
         \ML_int[4][3] , \ML_int[4][2] , n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14;
  assign B[11] = \ML_int[4][11] ;
  assign B[10] = \ML_int[4][10] ;
  assign B[9] = \ML_int[4][9] ;
  assign B[8] = \ML_int[4][8] ;
  assign B[7] = \ML_int[4][7] ;
  assign B[6] = \ML_int[4][6] ;
  assign B[5] = \ML_int[4][5] ;
  assign B[4] = \ML_int[4][4] ;
  assign B[3] = \ML_int[4][3] ;
  assign B[2] = \ML_int[4][2] ;

  MUX2D0BWP M1_2_8 ( .I0(\ML_int[2][8] ), .I1(\ML_int[2][4] ), .S(SH[2]), .Z(
        \ML_int[3][8] ) );
  MUX2D1BWP M1_3_8 ( .I0(\ML_int[3][8] ), .I1(\ML_int[3][0] ), .S(SH[3]), .Z(
        \ML_int[4][8] ) );
  MUX2D0BWP M1_2_9 ( .I0(\ML_int[2][9] ), .I1(\ML_int[2][5] ), .S(SH[2]), .Z(
        \ML_int[3][9] ) );
  MUX2D1BWP M1_3_9 ( .I0(\ML_int[3][9] ), .I1(\ML_int[3][1] ), .S(SH[3]), .Z(
        \ML_int[4][9] ) );
  MUX2D1BWP M1_3_10 ( .I0(\ML_int[3][10] ), .I1(n7), .S(SH[3]), .Z(
        \ML_int[4][10] ) );
  MUX2D1BWP M1_3_11 ( .I0(\ML_int[3][11] ), .I1(n6), .S(SH[3]), .Z(
        \ML_int[4][11] ) );
  MUX2D0BWP M1_0_4 ( .I0(A[4]), .I1(A[3]), .S(SH[0]), .Z(\ML_int[1][4] ) );
  MUX2D0BWP M1_0_3 ( .I0(A[3]), .I1(A[2]), .S(SH[0]), .Z(\ML_int[1][3] ) );
  MUX2D0BWP M1_1_3 ( .I0(\ML_int[1][3] ), .I1(\ML_int[1][1] ), .S(SH[1]), .Z(
        \ML_int[2][3] ) );
  MUX2D0BWP M1_1_4 ( .I0(\ML_int[1][4] ), .I1(\ML_int[1][2] ), .S(SH[1]), .Z(
        \ML_int[2][4] ) );
  MUX2D0BWP M1_1_5 ( .I0(\ML_int[1][5] ), .I1(\ML_int[1][3] ), .S(SH[1]), .Z(
        \ML_int[2][5] ) );
  MUX2D0BWP M1_1_6 ( .I0(\ML_int[1][6] ), .I1(\ML_int[1][4] ), .S(SH[1]), .Z(
        \ML_int[2][6] ) );
  MUX2D0BWP M1_0_10 ( .I0(A[10]), .I1(A[9]), .S(SH[0]), .Z(\ML_int[1][10] ) );
  MUX2D0BWP M1_1_10 ( .I0(\ML_int[1][10] ), .I1(\ML_int[1][8] ), .S(SH[1]), 
        .Z(\ML_int[2][10] ) );
  MUX2D0BWP M1_2_10 ( .I0(\ML_int[2][10] ), .I1(\ML_int[2][6] ), .S(SH[2]), 
        .Z(\ML_int[3][10] ) );
  MUX2D0BWP M1_0_11 ( .I0(A[11]), .I1(A[10]), .S(SH[0]), .Z(\ML_int[1][11] )
         );
  MUX2D0BWP M1_1_11 ( .I0(\ML_int[1][11] ), .I1(\ML_int[1][9] ), .S(SH[1]), 
        .Z(\ML_int[2][11] ) );
  MUX2D0BWP M1_2_11 ( .I0(\ML_int[2][11] ), .I1(\ML_int[2][7] ), .S(SH[2]), 
        .Z(\ML_int[3][11] ) );
  MUX2D0BWP M1_0_1 ( .I0(A[1]), .I1(A[0]), .S(SH[0]), .Z(\ML_int[1][1] ) );
  MUX2D0BWP M1_0_2 ( .I0(A[2]), .I1(A[1]), .S(SH[0]), .Z(\ML_int[1][2] ) );
  MUX2D0BWP M1_0_5 ( .I0(A[5]), .I1(A[4]), .S(SH[0]), .Z(\ML_int[1][5] ) );
  MUX2D0BWP M1_0_6 ( .I0(A[6]), .I1(A[5]), .S(SH[0]), .Z(\ML_int[1][6] ) );
  MUX2D0BWP M1_0_7 ( .I0(A[7]), .I1(A[6]), .S(SH[0]), .Z(\ML_int[1][7] ) );
  MUX2D0BWP M1_0_8 ( .I0(A[8]), .I1(A[7]), .S(SH[0]), .Z(\ML_int[1][8] ) );
  MUX2D0BWP M1_0_9 ( .I0(A[9]), .I1(A[8]), .S(SH[0]), .Z(\ML_int[1][9] ) );
  MUX2D0BWP M1_1_8 ( .I0(\ML_int[1][8] ), .I1(\ML_int[1][6] ), .S(SH[1]), .Z(
        \ML_int[2][8] ) );
  MUX2D0BWP M1_1_9 ( .I0(\ML_int[1][9] ), .I1(\ML_int[1][7] ), .S(SH[1]), .Z(
        \ML_int[2][9] ) );
  MUX2D0BWP M1_1_2 ( .I0(\ML_int[1][2] ), .I1(\ML_int[1][0] ), .S(SH[1]), .Z(
        \ML_int[2][2] ) );
  MUX2D0BWP M1_1_7 ( .I0(\ML_int[1][7] ), .I1(\ML_int[1][5] ), .S(SH[1]), .Z(
        \ML_int[2][7] ) );
  CKND0BWP U3 ( .I(SH[2]), .ZN(n9) );
  INVD1BWP U4 ( .I(SH[1]), .ZN(n10) );
  INVD1BWP U5 ( .I(n13), .ZN(n5) );
  INVD1BWP U6 ( .I(n14), .ZN(n8) );
  INR2D1BWP U7 ( .A1(A[0]), .B1(SH[0]), .ZN(\ML_int[1][0] ) );
  INVD1BWP U8 ( .I(n11), .ZN(n6) );
  INVD1BWP U9 ( .I(n12), .ZN(n7) );
  NR2XD0BWP U10 ( .A1(n1), .A2(SH[3]), .ZN(\ML_int[4][7] ) );
  MUX2ND0BWP U11 ( .I0(\ML_int[2][7] ), .I1(\ML_int[2][3] ), .S(SH[2]), .ZN(n1) );
  NR2XD0BWP U12 ( .A1(n2), .A2(SH[3]), .ZN(\ML_int[4][6] ) );
  MUX2ND0BWP U13 ( .I0(\ML_int[2][6] ), .I1(\ML_int[2][2] ), .S(SH[2]), .ZN(n2) );
  NR2XD0BWP U14 ( .A1(n3), .A2(SH[3]), .ZN(\ML_int[4][5] ) );
  MUX2ND0BWP U15 ( .I0(\ML_int[2][5] ), .I1(n5), .S(SH[2]), .ZN(n3) );
  NR2XD0BWP U16 ( .A1(n4), .A2(SH[3]), .ZN(\ML_int[4][4] ) );
  MUX2ND0BWP U17 ( .I0(\ML_int[2][4] ), .I1(n8), .S(SH[2]), .ZN(n4) );
  NR2D0BWP U18 ( .A1(n11), .A2(SH[3]), .ZN(\ML_int[4][3] ) );
  NR2D0BWP U19 ( .A1(n12), .A2(SH[3]), .ZN(\ML_int[4][2] ) );
  CKND2D0BWP U20 ( .A1(\ML_int[2][3] ), .A2(n9), .ZN(n11) );
  CKND2D0BWP U21 ( .A1(\ML_int[2][2] ), .A2(n9), .ZN(n12) );
  NR2D0BWP U22 ( .A1(SH[2]), .A2(n13), .ZN(\ML_int[3][1] ) );
  NR2D0BWP U23 ( .A1(SH[2]), .A2(n14), .ZN(\ML_int[3][0] ) );
  CKND2D0BWP U24 ( .A1(\ML_int[1][1] ), .A2(n10), .ZN(n13) );
  CKND2D0BWP U25 ( .A1(\ML_int[1][0] ), .A2(n10), .ZN(n14) );
endmodule


module CVP14_DW01_addsub_3 ( A, B, CI, ADD_SUB, SUM, CO );
  input [5:0] A;
  input [5:0] B;
  output [5:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [6:0] carry;
  wire   [5:0] B_AS;
  assign carry[0] = ADD_SUB;

  FA1D0BWP U1_4 ( .A(A[4]), .B(carry[0]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FA1D0BWP U1_0 ( .A(A[0]), .B(B_AS[0]), .CI(carry[0]), .CO(carry[1]), .S(
        SUM[0]) );
  XOR3D1BWP U1_5 ( .A1(A[5]), .A2(carry[0]), .A3(carry[5]), .Z(SUM[5]) );
  FA1D0BWP U1_1 ( .A(A[1]), .B(B_AS[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  FA1D0BWP U1_3 ( .A(A[3]), .B(B_AS[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FA1D0BWP U1_2 ( .A(A[2]), .B(B_AS[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  CKXOR2D0BWP U1 ( .A1(B[3]), .A2(carry[0]), .Z(B_AS[3]) );
  CKXOR2D0BWP U2 ( .A1(B[2]), .A2(carry[0]), .Z(B_AS[2]) );
  CKXOR2D0BWP U3 ( .A1(B[1]), .A2(carry[0]), .Z(B_AS[1]) );
  CKXOR2D0BWP U4 ( .A1(B[0]), .A2(carry[0]), .Z(B_AS[0]) );
endmodule


module CVP14_DW01_inc_2 ( A, SUM );
  input [26:0] A;
  output [26:0] SUM;
  wire   n1, n2, n3, n4;
  wire   [26:2] carry;

  HA1D0BWP U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  HA1D0BWP U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  HA1D0BWP U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(SUM[26]), .S(SUM[25]) );
  HA1D0BWP U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  HA1D0BWP U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  HA1D0BWP U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  HA1D0BWP U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  HA1D0BWP U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  HA1D0BWP U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  HA1D0BWP U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  HA1D0BWP U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  HA1D0BWP U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  HA1D0BWP U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  NR4D0BWP U1 ( .A1(n1), .A2(n2), .A3(n3), .A4(n4), .ZN(carry[13]) );
  ND3D0BWP U2 ( .A1(A[8]), .A2(A[7]), .A3(A[9]), .ZN(n4) );
  ND3D0BWP U3 ( .A1(A[5]), .A2(A[4]), .A3(A[6]), .ZN(n3) );
  ND3D0BWP U4 ( .A1(A[2]), .A2(A[1]), .A3(A[3]), .ZN(n2) );
  ND4D0BWP U5 ( .A1(A[12]), .A2(A[11]), .A3(A[10]), .A4(A[0]), .ZN(n1) );
endmodule


module CVP14_DW01_ash_5 ( A, DATA_TC, SH, SH_TC, B );
  input [12:0] A;
  input [3:0] SH;
  output [12:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][12] , \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] ,
         \ML_int[1][8] , \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] ,
         \ML_int[1][4] , \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] ,
         \ML_int[1][0] , \ML_int[2][12] , \ML_int[2][11] , \ML_int[2][10] ,
         \ML_int[2][9] , \ML_int[2][8] , \ML_int[2][7] , \ML_int[2][6] ,
         \ML_int[2][5] , \ML_int[2][4] , \ML_int[2][3] , \ML_int[2][2] ,
         \ML_int[3][12] , \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] ,
         \ML_int[3][8] , \ML_int[3][5] , \ML_int[3][4] , \ML_int[3][3] ,
         \ML_int[3][2] , \ML_int[3][1] , \ML_int[3][0] , \ML_int[4][12] ,
         \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] ,
         \ML_int[4][7] , \ML_int[4][6] , \ML_int[4][5] , \ML_int[4][4] ,
         \ML_int[4][3] , \ML_int[4][2] , \ML_int[4][1] , \ML_int[4][0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10;
  assign B[12] = \ML_int[4][12] ;
  assign B[11] = \ML_int[4][11] ;
  assign B[10] = \ML_int[4][10] ;
  assign B[9] = \ML_int[4][9] ;
  assign B[8] = \ML_int[4][8] ;
  assign B[7] = \ML_int[4][7] ;
  assign B[6] = \ML_int[4][6] ;
  assign B[5] = \ML_int[4][5] ;
  assign B[4] = \ML_int[4][4] ;
  assign B[3] = \ML_int[4][3] ;
  assign B[2] = \ML_int[4][2] ;
  assign B[1] = \ML_int[4][1] ;
  assign B[0] = \ML_int[4][0] ;

  MUX2D0BWP M1_0_4 ( .I0(A[4]), .I1(A[3]), .S(SH[0]), .Z(\ML_int[1][4] ) );
  MUX2D0BWP M1_0_3 ( .I0(A[3]), .I1(A[2]), .S(SH[0]), .Z(\ML_int[1][3] ) );
  MUX2D0BWP M1_0_11 ( .I0(A[11]), .I1(A[10]), .S(SH[0]), .Z(\ML_int[1][11] )
         );
  MUX2D0BWP M1_1_11 ( .I0(\ML_int[1][11] ), .I1(\ML_int[1][9] ), .S(SH[1]), 
        .Z(\ML_int[2][11] ) );
  MUX2D0BWP M1_1_6 ( .I0(\ML_int[1][6] ), .I1(\ML_int[1][4] ), .S(SH[1]), .Z(
        \ML_int[2][6] ) );
  MUX2D0BWP M1_1_5 ( .I0(\ML_int[1][5] ), .I1(\ML_int[1][3] ), .S(SH[1]), .Z(
        \ML_int[2][5] ) );
  MUX2D0BWP M1_1_4 ( .I0(\ML_int[1][4] ), .I1(\ML_int[1][2] ), .S(SH[1]), .Z(
        \ML_int[2][4] ) );
  MUX2D0BWP M1_0_12 ( .I0(A[12]), .I1(A[11]), .S(SH[0]), .Z(\ML_int[1][12] )
         );
  MUX2D0BWP M1_0_10 ( .I0(A[10]), .I1(A[9]), .S(SH[0]), .Z(\ML_int[1][10] ) );
  MUX2D0BWP M1_0_8 ( .I0(A[8]), .I1(A[7]), .S(SH[0]), .Z(\ML_int[1][8] ) );
  MUX2D0BWP M1_0_6 ( .I0(A[6]), .I1(A[5]), .S(SH[0]), .Z(\ML_int[1][6] ) );
  MUX2D0BWP M1_0_9 ( .I0(A[9]), .I1(A[8]), .S(SH[0]), .Z(\ML_int[1][9] ) );
  MUX2D0BWP M1_0_7 ( .I0(A[7]), .I1(A[6]), .S(SH[0]), .Z(\ML_int[1][7] ) );
  MUX2D0BWP M1_0_5 ( .I0(A[5]), .I1(A[4]), .S(SH[0]), .Z(\ML_int[1][5] ) );
  MUX2D0BWP M1_0_2 ( .I0(A[2]), .I1(A[1]), .S(SH[0]), .Z(\ML_int[1][2] ) );
  MUX2D0BWP M1_1_3 ( .I0(\ML_int[1][3] ), .I1(\ML_int[1][1] ), .S(SH[1]), .Z(
        \ML_int[2][3] ) );
  MUX2D0BWP M1_1_12 ( .I0(\ML_int[1][12] ), .I1(\ML_int[1][10] ), .S(SH[1]), 
        .Z(\ML_int[2][12] ) );
  MUX2D0BWP M1_2_12 ( .I0(\ML_int[2][12] ), .I1(\ML_int[2][8] ), .S(SH[2]), 
        .Z(\ML_int[3][12] ) );
  MUX2D1BWP M1_3_12 ( .I0(\ML_int[3][12] ), .I1(\ML_int[3][4] ), .S(SH[3]), 
        .Z(\ML_int[4][12] ) );
  MUX2D0BWP M1_2_10 ( .I0(\ML_int[2][10] ), .I1(\ML_int[2][6] ), .S(SH[2]), 
        .Z(\ML_int[3][10] ) );
  MUX2D1BWP M1_3_10 ( .I0(\ML_int[3][10] ), .I1(\ML_int[3][2] ), .S(SH[3]), 
        .Z(\ML_int[4][10] ) );
  MUX2D0BWP M1_2_9 ( .I0(\ML_int[2][9] ), .I1(\ML_int[2][5] ), .S(SH[2]), .Z(
        \ML_int[3][9] ) );
  MUX2D1BWP M1_3_9 ( .I0(\ML_int[3][9] ), .I1(\ML_int[3][1] ), .S(SH[3]), .Z(
        \ML_int[4][9] ) );
  MUX2D0BWP M1_2_5 ( .I0(\ML_int[2][5] ), .I1(n3), .S(SH[2]), .Z(
        \ML_int[3][5] ) );
  MUX2D0BWP M1_2_11 ( .I0(\ML_int[2][11] ), .I1(\ML_int[2][7] ), .S(SH[2]), 
        .Z(\ML_int[3][11] ) );
  MUX2D1BWP M1_3_11 ( .I0(\ML_int[3][11] ), .I1(\ML_int[3][3] ), .S(SH[3]), 
        .Z(\ML_int[4][11] ) );
  MUX2D0BWP M1_2_8 ( .I0(\ML_int[2][8] ), .I1(\ML_int[2][4] ), .S(SH[2]), .Z(
        \ML_int[3][8] ) );
  MUX2D1BWP M1_3_8 ( .I0(\ML_int[3][8] ), .I1(\ML_int[3][0] ), .S(SH[3]), .Z(
        \ML_int[4][8] ) );
  MUX2D0BWP M1_1_10 ( .I0(\ML_int[1][10] ), .I1(\ML_int[1][8] ), .S(SH[1]), 
        .Z(\ML_int[2][10] ) );
  MUX2D0BWP M1_1_9 ( .I0(\ML_int[1][9] ), .I1(\ML_int[1][7] ), .S(SH[1]), .Z(
        \ML_int[2][9] ) );
  MUX2D0BWP M1_1_8 ( .I0(\ML_int[1][8] ), .I1(\ML_int[1][6] ), .S(SH[1]), .Z(
        \ML_int[2][8] ) );
  MUX2D0BWP M1_1_7 ( .I0(\ML_int[1][7] ), .I1(\ML_int[1][5] ), .S(SH[1]), .Z(
        \ML_int[2][7] ) );
  MUX2D0BWP M1_0_1 ( .I0(A[1]), .I1(A[0]), .S(SH[0]), .Z(\ML_int[1][1] ) );
  MUX2D1BWP M1_1_2 ( .I0(\ML_int[1][2] ), .I1(\ML_int[1][0] ), .S(SH[1]), .Z(
        \ML_int[2][2] ) );
  MUX2D0BWP M1_2_4 ( .I0(\ML_int[2][4] ), .I1(n4), .S(SH[2]), .Z(
        \ML_int[3][4] ) );
  OR2D0BWP U3 ( .A1(SH[3]), .A2(SH[2]), .Z(n8) );
  INVD1BWP U4 ( .I(\ML_int[2][2] ), .ZN(n6) );
  INVD1BWP U5 ( .I(n10), .ZN(n4) );
  INVD1BWP U6 ( .I(SH[1]), .ZN(n5) );
  INVD1BWP U7 ( .I(\ML_int[2][3] ), .ZN(n7) );
  NR2XD0BWP U8 ( .A1(n1), .A2(SH[3]), .ZN(\ML_int[4][7] ) );
  MUX2ND0BWP U9 ( .I0(\ML_int[2][7] ), .I1(\ML_int[2][3] ), .S(SH[2]), .ZN(n1)
         );
  INVD1BWP U10 ( .I(n9), .ZN(n3) );
  NR2XD0BWP U11 ( .A1(n2), .A2(SH[3]), .ZN(\ML_int[4][6] ) );
  MUX2ND0BWP U12 ( .I0(\ML_int[2][6] ), .I1(\ML_int[2][2] ), .S(SH[2]), .ZN(n2) );
  INR2D0BWP U13 ( .A1(\ML_int[3][5] ), .B1(SH[3]), .ZN(\ML_int[4][5] ) );
  INR2D0BWP U14 ( .A1(\ML_int[3][4] ), .B1(SH[3]), .ZN(\ML_int[4][4] ) );
  NR2D0BWP U15 ( .A1(n8), .A2(n7), .ZN(\ML_int[4][3] ) );
  NR2D0BWP U16 ( .A1(n8), .A2(n6), .ZN(\ML_int[4][2] ) );
  NR2D0BWP U17 ( .A1(n8), .A2(n9), .ZN(\ML_int[4][1] ) );
  NR2D0BWP U18 ( .A1(n8), .A2(n10), .ZN(\ML_int[4][0] ) );
  NR2D0BWP U19 ( .A1(SH[2]), .A2(n7), .ZN(\ML_int[3][3] ) );
  NR2D0BWP U20 ( .A1(SH[2]), .A2(n6), .ZN(\ML_int[3][2] ) );
  NR2D0BWP U21 ( .A1(SH[2]), .A2(n9), .ZN(\ML_int[3][1] ) );
  NR2D0BWP U22 ( .A1(SH[2]), .A2(n10), .ZN(\ML_int[3][0] ) );
  CKND2D0BWP U23 ( .A1(\ML_int[1][1] ), .A2(n5), .ZN(n9) );
  CKND2D0BWP U24 ( .A1(\ML_int[1][0] ), .A2(n5), .ZN(n10) );
  INR2D0BWP U25 ( .A1(A[0]), .B1(SH[0]), .ZN(\ML_int[1][0] ) );
endmodule


module CVP14_DW01_addsub_5 ( A, B, CI, ADD_SUB, SUM, CO );
  input [4:0] A;
  input [4:0] B;
  output [4:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [5:0] carry;
  wire   [4:0] B_AS;
  assign carry[0] = ADD_SUB;

  FA1D0BWP U1_3 ( .A(A[3]), .B(B_AS[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FA1D0BWP U1_2 ( .A(A[2]), .B(B_AS[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FA1D0BWP U1_1 ( .A(A[1]), .B(B_AS[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  FA1D0BWP U1_0 ( .A(A[0]), .B(B_AS[0]), .CI(carry[0]), .CO(carry[1]), .S(
        SUM[0]) );
  XOR3D1BWP U1_4 ( .A1(A[4]), .A2(carry[0]), .A3(carry[4]), .Z(SUM[4]) );
  CKXOR2D0BWP U1 ( .A1(B[3]), .A2(carry[0]), .Z(B_AS[3]) );
  CKXOR2D0BWP U2 ( .A1(B[2]), .A2(carry[0]), .Z(B_AS[2]) );
  CKXOR2D0BWP U3 ( .A1(B[1]), .A2(carry[0]), .Z(B_AS[1]) );
  CKXOR2D0BWP U4 ( .A1(B[0]), .A2(carry[0]), .Z(B_AS[0]) );
endmodule


module CVP14_DW01_addsub_6 ( A, B, CI, ADD_SUB, SUM, CO );
  input [26:0] A;
  input [26:0] B;
  output [26:0] SUM;
  input CI, ADD_SUB;
  output CO;
  wire   n1, n2;
  wire   [27:0] carry;
  wire   [26:0] B_AS;
  assign carry[0] = ADD_SUB;

  FA1D0BWP U1_16 ( .A(A[16]), .B(B_AS[16]), .CI(carry[16]), .CO(carry[17]), 
        .S(SUM[16]) );
  FA1D0BWP U1_24 ( .A(A[24]), .B(B_AS[24]), .CI(carry[24]), .CO(carry[25]), 
        .S(SUM[24]) );
  FA1D0BWP U1_23 ( .A(A[23]), .B(B_AS[23]), .CI(carry[23]), .CO(carry[24]), 
        .S(SUM[23]) );
  FA1D0BWP U1_22 ( .A(A[22]), .B(B_AS[22]), .CI(carry[22]), .CO(carry[23]), 
        .S(SUM[22]) );
  FA1D0BWP U1_21 ( .A(A[21]), .B(B_AS[21]), .CI(carry[21]), .CO(carry[22]), 
        .S(SUM[21]) );
  FA1D0BWP U1_19 ( .A(A[19]), .B(B_AS[19]), .CI(carry[19]), .CO(carry[20]), 
        .S(SUM[19]) );
  FA1D0BWP U1_17 ( .A(A[17]), .B(B_AS[17]), .CI(carry[17]), .CO(carry[18]), 
        .S(SUM[17]) );
  FA1D0BWP U1_20 ( .A(A[20]), .B(B_AS[20]), .CI(carry[20]), .CO(carry[21]), 
        .S(SUM[20]) );
  FA1D0BWP U1_15 ( .A(A[15]), .B(B_AS[15]), .CI(carry[15]), .CO(carry[16]), 
        .S(SUM[15]) );
  FA1D0BWP U1_18 ( .A(A[18]), .B(B_AS[18]), .CI(carry[18]), .CO(carry[19]), 
        .S(SUM[18]) );
  FA1D0BWP U1_25 ( .A(A[25]), .B(B_AS[25]), .CI(carry[25]), .CO(carry[26]), 
        .S(SUM[25]) );
  INVD1BWP U1 ( .I(carry[14]), .ZN(n2) );
  INVD1BWP U2 ( .I(B_AS[14]), .ZN(n1) );
  XOR2D1BWP U3 ( .A1(carry[14]), .A2(B_AS[14]), .Z(SUM[14]) );
  AN2XD1BWP U4 ( .A1(B_AS[1]), .A2(carry[1]), .Z(carry[2]) );
  AN2XD1BWP U5 ( .A1(B_AS[2]), .A2(carry[2]), .Z(carry[3]) );
  AN2XD1BWP U6 ( .A1(B_AS[3]), .A2(carry[3]), .Z(carry[4]) );
  AN2XD1BWP U7 ( .A1(B_AS[4]), .A2(carry[4]), .Z(carry[5]) );
  AN2XD1BWP U8 ( .A1(B_AS[5]), .A2(carry[5]), .Z(carry[6]) );
  AN2XD1BWP U9 ( .A1(B_AS[6]), .A2(carry[6]), .Z(carry[7]) );
  AN2XD1BWP U10 ( .A1(B_AS[7]), .A2(carry[7]), .Z(carry[8]) );
  AN2XD1BWP U11 ( .A1(B_AS[8]), .A2(carry[8]), .Z(carry[9]) );
  AN2XD1BWP U12 ( .A1(B_AS[9]), .A2(carry[9]), .Z(carry[10]) );
  AN2XD1BWP U13 ( .A1(B_AS[10]), .A2(carry[10]), .Z(carry[11]) );
  AN2XD1BWP U14 ( .A1(B_AS[11]), .A2(carry[11]), .Z(carry[12]) );
  AN2XD1BWP U15 ( .A1(B_AS[12]), .A2(carry[12]), .Z(carry[13]) );
  AN2XD1BWP U16 ( .A1(B_AS[13]), .A2(carry[13]), .Z(carry[14]) );
  XOR2D1BWP U17 ( .A1(carry[13]), .A2(B_AS[13]), .Z(SUM[13]) );
  XOR2D1BWP U18 ( .A1(carry[5]), .A2(B_AS[5]), .Z(SUM[5]) );
  XOR2D1BWP U19 ( .A1(carry[9]), .A2(B_AS[9]), .Z(SUM[9]) );
  XOR2D1BWP U20 ( .A1(carry[1]), .A2(B_AS[1]), .Z(SUM[1]) );
  XOR2D1BWP U21 ( .A1(carry[6]), .A2(B_AS[6]), .Z(SUM[6]) );
  XOR2D1BWP U22 ( .A1(carry[10]), .A2(B_AS[10]), .Z(SUM[10]) );
  XOR2D1BWP U23 ( .A1(carry[2]), .A2(B_AS[2]), .Z(SUM[2]) );
  XOR2D1BWP U24 ( .A1(carry[7]), .A2(B_AS[7]), .Z(SUM[7]) );
  XOR2D1BWP U25 ( .A1(carry[11]), .A2(B_AS[11]), .Z(SUM[11]) );
  XOR2D1BWP U26 ( .A1(carry[3]), .A2(B_AS[3]), .Z(SUM[3]) );
  XOR2D1BWP U27 ( .A1(carry[8]), .A2(B_AS[8]), .Z(SUM[8]) );
  XOR2D1BWP U28 ( .A1(carry[12]), .A2(B_AS[12]), .Z(SUM[12]) );
  XOR2D1BWP U29 ( .A1(carry[4]), .A2(B_AS[4]), .Z(SUM[4]) );
  XOR2D1BWP U30 ( .A1(carry[0]), .A2(carry[26]), .Z(SUM[26]) );
  AN2XD1BWP U31 ( .A1(B_AS[0]), .A2(carry[0]), .Z(carry[1]) );
  CKXOR2D0BWP U32 ( .A1(carry[0]), .A2(B_AS[0]), .Z(SUM[0]) );
  NR2XD0BWP U33 ( .A1(n1), .A2(n2), .ZN(carry[15]) );
  CKXOR2D0BWP U34 ( .A1(B[9]), .A2(carry[0]), .Z(B_AS[9]) );
  CKXOR2D0BWP U35 ( .A1(B[8]), .A2(carry[0]), .Z(B_AS[8]) );
  CKXOR2D0BWP U36 ( .A1(B[7]), .A2(carry[0]), .Z(B_AS[7]) );
  CKXOR2D0BWP U37 ( .A1(B[6]), .A2(carry[0]), .Z(B_AS[6]) );
  CKXOR2D0BWP U38 ( .A1(B[5]), .A2(carry[0]), .Z(B_AS[5]) );
  CKXOR2D0BWP U39 ( .A1(B[4]), .A2(carry[0]), .Z(B_AS[4]) );
  CKXOR2D0BWP U40 ( .A1(B[3]), .A2(carry[0]), .Z(B_AS[3]) );
  CKXOR2D0BWP U41 ( .A1(B[2]), .A2(carry[0]), .Z(B_AS[2]) );
  CKXOR2D0BWP U42 ( .A1(B[25]), .A2(carry[0]), .Z(B_AS[25]) );
  CKXOR2D0BWP U43 ( .A1(B[24]), .A2(carry[0]), .Z(B_AS[24]) );
  CKXOR2D0BWP U44 ( .A1(B[23]), .A2(carry[0]), .Z(B_AS[23]) );
  CKXOR2D0BWP U45 ( .A1(B[22]), .A2(carry[0]), .Z(B_AS[22]) );
  CKXOR2D0BWP U46 ( .A1(B[21]), .A2(carry[0]), .Z(B_AS[21]) );
  CKXOR2D0BWP U47 ( .A1(B[20]), .A2(carry[0]), .Z(B_AS[20]) );
  CKXOR2D0BWP U48 ( .A1(B[1]), .A2(carry[0]), .Z(B_AS[1]) );
  CKXOR2D0BWP U49 ( .A1(B[19]), .A2(carry[0]), .Z(B_AS[19]) );
  CKXOR2D0BWP U50 ( .A1(B[18]), .A2(carry[0]), .Z(B_AS[18]) );
  CKXOR2D0BWP U51 ( .A1(B[17]), .A2(carry[0]), .Z(B_AS[17]) );
  CKXOR2D0BWP U52 ( .A1(B[16]), .A2(carry[0]), .Z(B_AS[16]) );
  CKXOR2D0BWP U53 ( .A1(B[15]), .A2(carry[0]), .Z(B_AS[15]) );
  CKXOR2D0BWP U54 ( .A1(B[14]), .A2(carry[0]), .Z(B_AS[14]) );
  CKXOR2D0BWP U55 ( .A1(B[13]), .A2(carry[0]), .Z(B_AS[13]) );
  CKXOR2D0BWP U56 ( .A1(B[12]), .A2(carry[0]), .Z(B_AS[12]) );
  CKXOR2D0BWP U57 ( .A1(B[11]), .A2(carry[0]), .Z(B_AS[11]) );
  CKXOR2D0BWP U58 ( .A1(B[10]), .A2(carry[0]), .Z(B_AS[10]) );
  CKXOR2D0BWP U59 ( .A1(B[0]), .A2(carry[0]), .Z(B_AS[0]) );
endmodule


module CVP14_DW_rash_2 ( A, DATA_TC, SH, SH_TC, B );
  input [25:0] A;
  input [4:0] SH;
  output [25:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76;

  INVD1BWP U3 ( .I(n65), .ZN(n16) );
  INVD1BWP U4 ( .I(n36), .ZN(n1) );
  INVD1BWP U5 ( .I(n34), .ZN(n4) );
  INVD1BWP U6 ( .I(n66), .ZN(n11) );
  INVD1BWP U7 ( .I(n58), .ZN(n6) );
  INVD1BWP U8 ( .I(n57), .ZN(n7) );
  INVD1BWP U9 ( .I(n67), .ZN(n2) );
  INVD1BWP U10 ( .I(n52), .ZN(n3) );
  INVD1BWP U11 ( .I(n41), .ZN(n10) );
  INVD1BWP U12 ( .I(n37), .ZN(n14) );
  INVD1BWP U13 ( .I(n40), .ZN(n15) );
  INVD1BWP U14 ( .I(SH[4]), .ZN(n5) );
  INVD1BWP U15 ( .I(SH[2]), .ZN(n8) );
  INVD1BWP U16 ( .I(SH[1]), .ZN(n17) );
  INVD1BWP U17 ( .I(SH[0]), .ZN(n18) );
  INVD1BWP U18 ( .I(A[25]), .ZN(n19) );
  INVD1BWP U19 ( .I(n56), .ZN(n12) );
  INVD1BWP U20 ( .I(n38), .ZN(n13) );
  INVD1BWP U21 ( .I(n69), .ZN(n9) );
  INVD1BWP U22 ( .I(A[17]), .ZN(n27) );
  INVD1BWP U23 ( .I(A[22]), .ZN(n22) );
  INVD1BWP U24 ( .I(A[21]), .ZN(n23) );
  INVD1BWP U25 ( .I(A[20]), .ZN(n24) );
  INVD1BWP U26 ( .I(A[19]), .ZN(n25) );
  INVD1BWP U27 ( .I(A[18]), .ZN(n26) );
  INVD1BWP U28 ( .I(A[15]), .ZN(n29) );
  INVD1BWP U29 ( .I(A[16]), .ZN(n28) );
  INVD1BWP U30 ( .I(A[24]), .ZN(n20) );
  INVD1BWP U31 ( .I(A[23]), .ZN(n21) );
  OAI221D0BWP U32 ( .A1(n30), .A2(n31), .B1(n13), .B2(n32), .C(n33), .ZN(B[9])
         );
  AOI22D0BWP U33 ( .A1(n34), .A2(n35), .B1(n36), .B2(n37), .ZN(n33) );
  OAI221D0BWP U34 ( .A1(n9), .A2(n31), .B1(n12), .B2(n32), .C(n39), .ZN(B[8])
         );
  AOI22D0BWP U35 ( .A1(n40), .A2(n36), .B1(n34), .B2(n41), .ZN(n39) );
  OAI222D0BWP U36 ( .A1(n42), .A2(n31), .B1(n43), .B2(n4), .C1(n44), .C2(n32), 
        .ZN(B[7]) );
  OAI222D0BWP U37 ( .A1(n45), .A2(n31), .B1(n46), .B2(n4), .C1(n47), .C2(n32), 
        .ZN(B[6]) );
  NR2D0BWP U38 ( .A1(n5), .A2(n7), .ZN(n34) );
  OAI21D0BWP U39 ( .A1(n30), .A2(n32), .B(n48), .ZN(B[5]) );
  OA32D0BWP U40 ( .A1(n49), .A2(SH[3]), .A3(n5), .B1(n31), .B2(n14), .Z(n48)
         );
  OAI22D0BWP U41 ( .A1(n50), .A2(n5), .B1(n51), .B2(n52), .ZN(B[4]) );
  OAI22D0BWP U42 ( .A1(n53), .A2(n5), .B1(n42), .B2(n32), .ZN(B[3]) );
  OAI22D0BWP U43 ( .A1(n54), .A2(n5), .B1(n45), .B2(n32), .ZN(B[2]) );
  INR2D0BWP U44 ( .A1(n35), .B1(n55), .ZN(B[25]) );
  NR2D0BWP U45 ( .A1(n10), .A2(n55), .ZN(B[24]) );
  NR2D0BWP U46 ( .A1(n43), .A2(n55), .ZN(B[23]) );
  NR2D0BWP U47 ( .A1(n46), .A2(n55), .ZN(B[22]) );
  NR2D0BWP U48 ( .A1(n49), .A2(n2), .ZN(B[21]) );
  NR2D0BWP U49 ( .A1(SH[4]), .A2(n50), .ZN(B[20]) );
  AOI22D0BWP U50 ( .A1(n56), .A2(n57), .B1(n41), .B2(n58), .ZN(n50) );
  OAI22D0BWP U51 ( .A1(n59), .A2(n5), .B1(n14), .B2(n32), .ZN(B[1]) );
  NR2D0BWP U52 ( .A1(SH[4]), .A2(n53), .ZN(B[19]) );
  OA22D1BWP U53 ( .A1(n44), .A2(n7), .B1(n43), .B2(n6), .Z(n53) );
  NR2D0BWP U54 ( .A1(SH[4]), .A2(n54), .ZN(B[18]) );
  OA22D1BWP U55 ( .A1(n47), .A2(n7), .B1(n46), .B2(n6), .Z(n54) );
  NR2D0BWP U56 ( .A1(SH[4]), .A2(n59), .ZN(B[17]) );
  OA21D0BWP U57 ( .A1(n30), .A2(n7), .B(n60), .Z(n59) );
  AOI32D0BWP U58 ( .A1(n35), .A2(n8), .A3(SH[3]), .B1(n58), .B2(n38), .ZN(n60)
         );
  NR2D0BWP U59 ( .A1(SH[4]), .A2(n61), .ZN(B[16]) );
  OAI222D0BWP U60 ( .A1(n44), .A2(n1), .B1(n42), .B2(n55), .C1(n43), .C2(n31), 
        .ZN(B[15]) );
  OAI222D0BWP U61 ( .A1(n47), .A2(n1), .B1(n45), .B2(n55), .C1(n46), .C2(n31), 
        .ZN(B[14]) );
  OAI222D0BWP U62 ( .A1(n30), .A2(n1), .B1(n14), .B2(n55), .C1(n49), .C2(n52), 
        .ZN(B[13]) );
  MUX2ND0BWP U63 ( .I0(n35), .I1(n38), .S(n8), .ZN(n49) );
  OAI221D0BWP U64 ( .A1(n62), .A2(n22), .B1(n63), .B2(n21), .C(n64), .ZN(n38)
         );
  AOI22D0BWP U65 ( .A1(A[24]), .A2(n65), .B1(A[21]), .B2(n66), .ZN(n64) );
  NR2D0BWP U66 ( .A1(n19), .A2(n11), .ZN(n35) );
  CKND2D0BWP U67 ( .A1(n67), .A2(n8), .ZN(n55) );
  OAI22D0BWP U68 ( .A1(n16), .A2(n28), .B1(n63), .B2(n29), .ZN(n37) );
  OA221D0BWP U69 ( .A1(n62), .A2(n26), .B1(n63), .B2(n25), .C(n68), .Z(n30) );
  AOI22D0BWP U70 ( .A1(A[20]), .A2(n65), .B1(A[17]), .B2(n66), .ZN(n68) );
  OAI222D0BWP U71 ( .A1(n10), .A2(n32), .B1(n12), .B2(n31), .C1(n51), .C2(n2), 
        .ZN(B[12]) );
  MUX2ND0BWP U72 ( .I0(n69), .I1(n40), .S(n8), .ZN(n51) );
  OAI222D0BWP U73 ( .A1(n44), .A2(n31), .B1(n42), .B2(n1), .C1(n43), .C2(n32), 
        .ZN(B[11]) );
  OA222D0BWP U74 ( .A1(n19), .A2(n63), .B1(n62), .B2(n20), .C1(n11), .C2(n21), 
        .Z(n43) );
  OA221D0BWP U75 ( .A1(n28), .A2(n62), .B1(n63), .B2(n27), .C(n70), .Z(n42) );
  AOI22D0BWP U76 ( .A1(A[18]), .A2(n65), .B1(A[15]), .B2(n66), .ZN(n70) );
  OA221D0BWP U77 ( .A1(n62), .A2(n24), .B1(n63), .B2(n23), .C(n71), .Z(n44) );
  AOI22D0BWP U78 ( .A1(A[22]), .A2(n65), .B1(A[19]), .B2(n66), .ZN(n71) );
  OAI222D0BWP U79 ( .A1(n47), .A2(n31), .B1(n45), .B2(n1), .C1(n46), .C2(n32), 
        .ZN(B[10]) );
  OA221D0BWP U80 ( .A1(n62), .A2(n21), .B1(n63), .B2(n20), .C(n72), .Z(n46) );
  AOI22D0BWP U81 ( .A1(n65), .A2(A[25]), .B1(A[22]), .B2(n66), .ZN(n72) );
  NR2D0BWP U82 ( .A1(n8), .A2(n2), .ZN(n36) );
  NR2D0BWP U83 ( .A1(SH[3]), .A2(SH[4]), .ZN(n67) );
  OA222D0BWP U84 ( .A1(n63), .A2(n28), .B1(n29), .B2(n62), .C1(n16), .C2(n27), 
        .Z(n45) );
  CKND2D0BWP U85 ( .A1(n3), .A2(n8), .ZN(n31) );
  OA221D0BWP U86 ( .A1(n62), .A2(n25), .B1(n63), .B2(n24), .C(n73), .Z(n47) );
  AOI22D0BWP U87 ( .A1(A[21]), .A2(n65), .B1(A[18]), .B2(n66), .ZN(n73) );
  OAI22D0BWP U88 ( .A1(n61), .A2(n5), .B1(n32), .B2(n15), .ZN(B[0]) );
  NR2D0BWP U89 ( .A1(n16), .A2(n29), .ZN(n40) );
  CKND2D0BWP U90 ( .A1(n3), .A2(SH[2]), .ZN(n32) );
  CKND2D0BWP U91 ( .A1(SH[3]), .A2(n5), .ZN(n52) );
  OA21D0BWP U92 ( .A1(n9), .A2(n7), .B(n74), .Z(n61) );
  AOI32D0BWP U93 ( .A1(n41), .A2(n8), .A3(SH[3]), .B1(n58), .B2(n56), .ZN(n74)
         );
  OAI221D0BWP U94 ( .A1(n62), .A2(n23), .B1(n63), .B2(n22), .C(n75), .ZN(n56)
         );
  AOI22D0BWP U95 ( .A1(A[23]), .A2(n65), .B1(A[20]), .B2(n66), .ZN(n75) );
  NR2D0BWP U96 ( .A1(n8), .A2(SH[3]), .ZN(n58) );
  OAI22D0BWP U97 ( .A1(n11), .A2(n20), .B1(n19), .B2(n62), .ZN(n41) );
  NR2D0BWP U98 ( .A1(SH[2]), .A2(SH[3]), .ZN(n57) );
  OAI221D0BWP U99 ( .A1(n62), .A2(n27), .B1(n63), .B2(n26), .C(n76), .ZN(n69)
         );
  AOI22D0BWP U100 ( .A1(A[19]), .A2(n65), .B1(A[16]), .B2(n66), .ZN(n76) );
  NR2D0BWP U101 ( .A1(SH[0]), .A2(SH[1]), .ZN(n66) );
  NR2D0BWP U102 ( .A1(n18), .A2(n17), .ZN(n65) );
  CKND2D0BWP U103 ( .A1(SH[1]), .A2(n18), .ZN(n63) );
  CKND2D0BWP U104 ( .A1(SH[0]), .A2(n17), .ZN(n62) );
endmodule


module CVP14_DW_rash_3 ( A, DATA_TC, SH, SH_TC, B );
  input [25:0] A;
  input [4:0] SH;
  output [25:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76;

  INVD1BWP U3 ( .I(n65), .ZN(n16) );
  INVD1BWP U4 ( .I(n36), .ZN(n1) );
  INVD1BWP U5 ( .I(n34), .ZN(n4) );
  INVD1BWP U6 ( .I(n66), .ZN(n11) );
  INVD1BWP U7 ( .I(n58), .ZN(n6) );
  INVD1BWP U8 ( .I(n57), .ZN(n7) );
  INVD1BWP U9 ( .I(n67), .ZN(n2) );
  INVD1BWP U10 ( .I(n52), .ZN(n3) );
  INVD1BWP U11 ( .I(n41), .ZN(n10) );
  INVD1BWP U12 ( .I(n37), .ZN(n14) );
  INVD1BWP U13 ( .I(n40), .ZN(n15) );
  INVD1BWP U14 ( .I(SH[4]), .ZN(n5) );
  INVD1BWP U15 ( .I(SH[2]), .ZN(n8) );
  INVD1BWP U16 ( .I(SH[1]), .ZN(n17) );
  INVD1BWP U17 ( .I(SH[0]), .ZN(n18) );
  INVD1BWP U18 ( .I(A[25]), .ZN(n28) );
  INVD1BWP U19 ( .I(n56), .ZN(n12) );
  INVD1BWP U20 ( .I(n38), .ZN(n13) );
  INVD1BWP U21 ( .I(n69), .ZN(n9) );
  INVD1BWP U22 ( .I(A[15]), .ZN(n29) );
  INVD1BWP U23 ( .I(A[17]), .ZN(n21) );
  INVD1BWP U24 ( .I(A[21]), .ZN(n24) );
  INVD1BWP U25 ( .I(A[20]), .ZN(n23) );
  INVD1BWP U26 ( .I(A[19]), .ZN(n19) );
  INVD1BWP U27 ( .I(A[18]), .ZN(n20) );
  INVD1BWP U28 ( .I(A[16]), .ZN(n22) );
  INVD1BWP U29 ( .I(A[22]), .ZN(n25) );
  INVD1BWP U30 ( .I(A[24]), .ZN(n27) );
  INVD1BWP U31 ( .I(A[23]), .ZN(n26) );
  OAI221D0BWP U32 ( .A1(n30), .A2(n31), .B1(n13), .B2(n32), .C(n33), .ZN(B[9])
         );
  AOI22D0BWP U33 ( .A1(n34), .A2(n35), .B1(n36), .B2(n37), .ZN(n33) );
  OAI221D0BWP U34 ( .A1(n9), .A2(n31), .B1(n12), .B2(n32), .C(n39), .ZN(B[8])
         );
  AOI22D0BWP U35 ( .A1(n40), .A2(n36), .B1(n34), .B2(n41), .ZN(n39) );
  OAI222D0BWP U36 ( .A1(n42), .A2(n31), .B1(n43), .B2(n4), .C1(n44), .C2(n32), 
        .ZN(B[7]) );
  OAI222D0BWP U37 ( .A1(n45), .A2(n31), .B1(n46), .B2(n4), .C1(n47), .C2(n32), 
        .ZN(B[6]) );
  NR2D0BWP U38 ( .A1(n5), .A2(n7), .ZN(n34) );
  OAI21D0BWP U39 ( .A1(n30), .A2(n32), .B(n48), .ZN(B[5]) );
  OA32D0BWP U40 ( .A1(n49), .A2(SH[3]), .A3(n5), .B1(n31), .B2(n14), .Z(n48)
         );
  OAI22D0BWP U41 ( .A1(n50), .A2(n5), .B1(n51), .B2(n52), .ZN(B[4]) );
  OAI22D0BWP U42 ( .A1(n53), .A2(n5), .B1(n42), .B2(n32), .ZN(B[3]) );
  OAI22D0BWP U43 ( .A1(n54), .A2(n5), .B1(n45), .B2(n32), .ZN(B[2]) );
  INR2D0BWP U44 ( .A1(n35), .B1(n55), .ZN(B[25]) );
  NR2D0BWP U45 ( .A1(n10), .A2(n55), .ZN(B[24]) );
  NR2D0BWP U46 ( .A1(n43), .A2(n55), .ZN(B[23]) );
  NR2D0BWP U47 ( .A1(n46), .A2(n55), .ZN(B[22]) );
  NR2D0BWP U48 ( .A1(n49), .A2(n2), .ZN(B[21]) );
  NR2D0BWP U49 ( .A1(SH[4]), .A2(n50), .ZN(B[20]) );
  AOI22D0BWP U50 ( .A1(n56), .A2(n57), .B1(n41), .B2(n58), .ZN(n50) );
  OAI22D0BWP U51 ( .A1(n59), .A2(n5), .B1(n14), .B2(n32), .ZN(B[1]) );
  NR2D0BWP U52 ( .A1(SH[4]), .A2(n53), .ZN(B[19]) );
  OA22D1BWP U53 ( .A1(n44), .A2(n7), .B1(n43), .B2(n6), .Z(n53) );
  NR2D0BWP U54 ( .A1(SH[4]), .A2(n54), .ZN(B[18]) );
  OA22D1BWP U55 ( .A1(n47), .A2(n7), .B1(n46), .B2(n6), .Z(n54) );
  NR2D0BWP U56 ( .A1(SH[4]), .A2(n59), .ZN(B[17]) );
  OA21D0BWP U57 ( .A1(n30), .A2(n7), .B(n60), .Z(n59) );
  AOI32D0BWP U58 ( .A1(n35), .A2(n8), .A3(SH[3]), .B1(n58), .B2(n38), .ZN(n60)
         );
  NR2D0BWP U59 ( .A1(SH[4]), .A2(n61), .ZN(B[16]) );
  OAI222D0BWP U60 ( .A1(n44), .A2(n1), .B1(n42), .B2(n55), .C1(n43), .C2(n31), 
        .ZN(B[15]) );
  OAI222D0BWP U61 ( .A1(n47), .A2(n1), .B1(n45), .B2(n55), .C1(n46), .C2(n31), 
        .ZN(B[14]) );
  OAI222D0BWP U62 ( .A1(n30), .A2(n1), .B1(n14), .B2(n55), .C1(n49), .C2(n52), 
        .ZN(B[13]) );
  MUX2ND0BWP U63 ( .I0(n35), .I1(n38), .S(n8), .ZN(n49) );
  OAI221D0BWP U64 ( .A1(n62), .A2(n25), .B1(n63), .B2(n26), .C(n64), .ZN(n38)
         );
  AOI22D0BWP U65 ( .A1(A[24]), .A2(n65), .B1(A[21]), .B2(n66), .ZN(n64) );
  NR2D0BWP U66 ( .A1(n28), .A2(n11), .ZN(n35) );
  CKND2D0BWP U67 ( .A1(n67), .A2(n8), .ZN(n55) );
  OAI22D0BWP U68 ( .A1(n16), .A2(n22), .B1(n63), .B2(n29), .ZN(n37) );
  OA221D0BWP U69 ( .A1(n62), .A2(n20), .B1(n63), .B2(n19), .C(n68), .Z(n30) );
  AOI22D0BWP U70 ( .A1(A[20]), .A2(n65), .B1(A[17]), .B2(n66), .ZN(n68) );
  OAI222D0BWP U71 ( .A1(n10), .A2(n32), .B1(n12), .B2(n31), .C1(n51), .C2(n2), 
        .ZN(B[12]) );
  MUX2ND0BWP U72 ( .I0(n69), .I1(n40), .S(n8), .ZN(n51) );
  OAI222D0BWP U73 ( .A1(n44), .A2(n31), .B1(n42), .B2(n1), .C1(n43), .C2(n32), 
        .ZN(B[11]) );
  OA222D0BWP U74 ( .A1(n28), .A2(n63), .B1(n62), .B2(n27), .C1(n11), .C2(n26), 
        .Z(n43) );
  OA221D0BWP U75 ( .A1(n22), .A2(n62), .B1(n63), .B2(n21), .C(n70), .Z(n42) );
  AOI22D0BWP U76 ( .A1(A[18]), .A2(n65), .B1(A[15]), .B2(n66), .ZN(n70) );
  OA221D0BWP U77 ( .A1(n62), .A2(n23), .B1(n63), .B2(n24), .C(n71), .Z(n44) );
  AOI22D0BWP U78 ( .A1(A[22]), .A2(n65), .B1(A[19]), .B2(n66), .ZN(n71) );
  OAI222D0BWP U79 ( .A1(n47), .A2(n31), .B1(n45), .B2(n1), .C1(n46), .C2(n32), 
        .ZN(B[10]) );
  OA221D0BWP U80 ( .A1(n62), .A2(n26), .B1(n63), .B2(n27), .C(n72), .Z(n46) );
  AOI22D0BWP U81 ( .A1(n65), .A2(A[25]), .B1(A[22]), .B2(n66), .ZN(n72) );
  NR2D0BWP U82 ( .A1(n8), .A2(n2), .ZN(n36) );
  NR2D0BWP U83 ( .A1(SH[3]), .A2(SH[4]), .ZN(n67) );
  OA222D0BWP U84 ( .A1(n63), .A2(n22), .B1(n29), .B2(n62), .C1(n16), .C2(n21), 
        .Z(n45) );
  CKND2D0BWP U85 ( .A1(n3), .A2(n8), .ZN(n31) );
  OA221D0BWP U86 ( .A1(n62), .A2(n19), .B1(n63), .B2(n23), .C(n73), .Z(n47) );
  AOI22D0BWP U87 ( .A1(A[21]), .A2(n65), .B1(A[18]), .B2(n66), .ZN(n73) );
  OAI22D0BWP U88 ( .A1(n61), .A2(n5), .B1(n32), .B2(n15), .ZN(B[0]) );
  NR2D0BWP U89 ( .A1(n16), .A2(n29), .ZN(n40) );
  CKND2D0BWP U90 ( .A1(n3), .A2(SH[2]), .ZN(n32) );
  CKND2D0BWP U91 ( .A1(SH[3]), .A2(n5), .ZN(n52) );
  OA21D0BWP U92 ( .A1(n9), .A2(n7), .B(n74), .Z(n61) );
  AOI32D0BWP U93 ( .A1(n41), .A2(n8), .A3(SH[3]), .B1(n58), .B2(n56), .ZN(n74)
         );
  OAI221D0BWP U94 ( .A1(n62), .A2(n24), .B1(n63), .B2(n25), .C(n75), .ZN(n56)
         );
  AOI22D0BWP U95 ( .A1(A[23]), .A2(n65), .B1(A[20]), .B2(n66), .ZN(n75) );
  NR2D0BWP U96 ( .A1(n8), .A2(SH[3]), .ZN(n58) );
  OAI22D0BWP U97 ( .A1(n11), .A2(n27), .B1(n28), .B2(n62), .ZN(n41) );
  NR2D0BWP U98 ( .A1(SH[2]), .A2(SH[3]), .ZN(n57) );
  OAI221D0BWP U99 ( .A1(n62), .A2(n21), .B1(n63), .B2(n20), .C(n76), .ZN(n69)
         );
  AOI22D0BWP U100 ( .A1(A[19]), .A2(n65), .B1(A[16]), .B2(n66), .ZN(n76) );
  NR2D0BWP U101 ( .A1(SH[0]), .A2(SH[1]), .ZN(n66) );
  NR2D0BWP U102 ( .A1(n18), .A2(n17), .ZN(n65) );
  CKND2D0BWP U103 ( .A1(SH[1]), .A2(n18), .ZN(n63) );
  CKND2D0BWP U104 ( .A1(SH[0]), .A2(n17), .ZN(n62) );
endmodule


module CVP14_DW01_addsub_7 ( A, B, CI, ADD_SUB, SUM, CO );
  input [5:0] A;
  input [5:0] B;
  output [5:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [6:0] carry;
  wire   [5:0] B_AS;
  assign B_AS[5] = ADD_SUB;

  FA1D0BWP U1_0 ( .A(A[0]), .B(B_AS[0]), .CI(carry[0]), .CO(carry[1]), .S(
        SUM[0]) );
  FA1D0BWP U1_1 ( .A(A[1]), .B(B_AS[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  FA1D0BWP U1_3 ( .A(A[3]), .B(B_AS[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FA1D0BWP U1_4 ( .A(A[4]), .B(B_AS[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FA1D0BWP U1_2 ( .A(A[2]), .B(B_AS[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  XOR2D1BWP U1 ( .A1(B_AS[5]), .A2(carry[5]), .Z(SUM[5]) );
  CKXOR2D0BWP U2 ( .A1(CI), .A2(B_AS[5]), .Z(carry[0]) );
  CKXOR2D0BWP U3 ( .A1(B[4]), .A2(B_AS[5]), .Z(B_AS[4]) );
  CKXOR2D0BWP U4 ( .A1(B[3]), .A2(B_AS[5]), .Z(B_AS[3]) );
  CKXOR2D0BWP U5 ( .A1(B[2]), .A2(B_AS[5]), .Z(B_AS[2]) );
  CKXOR2D0BWP U6 ( .A1(B[1]), .A2(B_AS[5]), .Z(B_AS[1]) );
  CKXOR2D0BWP U7 ( .A1(B[0]), .A2(B_AS[5]), .Z(B_AS[0]) );
endmodule


module CVP14_DW01_decode_2 ( A, B );
  input [4:0] A;
  output [31:0] B;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;

  INVD1BWP U2 ( .I(A[2]), .ZN(n3) );
  INVD1BWP U3 ( .I(A[0]), .ZN(n2) );
  INVD1BWP U4 ( .I(A[3]), .ZN(n1) );
  NR2D0BWP U5 ( .A1(n4), .A2(n5), .ZN(B[9]) );
  NR2D0BWP U6 ( .A1(n4), .A2(n6), .ZN(B[8]) );
  NR2D0BWP U7 ( .A1(n7), .A2(n8), .ZN(B[7]) );
  NR2D0BWP U8 ( .A1(n7), .A2(n9), .ZN(B[6]) );
  NR2D0BWP U9 ( .A1(n8), .A2(n10), .ZN(B[5]) );
  NR2D0BWP U10 ( .A1(n9), .A2(n10), .ZN(B[4]) );
  NR2D0BWP U11 ( .A1(n8), .A2(n11), .ZN(B[3]) );
  NR2D0BWP U12 ( .A1(n9), .A2(n11), .ZN(B[2]) );
  NR2D0BWP U13 ( .A1(n4), .A2(n8), .ZN(B[1]) );
  CKND2D0BWP U14 ( .A1(A[0]), .A2(n1), .ZN(n8) );
  NR2D0BWP U15 ( .A1(n6), .A2(n7), .ZN(B[14]) );
  CKND2D0BWP U16 ( .A1(A[1]), .A2(n12), .ZN(n7) );
  NR2D0BWP U17 ( .A1(n5), .A2(n10), .ZN(B[13]) );
  NR2D0BWP U18 ( .A1(n6), .A2(n10), .ZN(B[12]) );
  IND2D0BWP U19 ( .A1(A[1]), .B1(n12), .ZN(n10) );
  NR2D0BWP U20 ( .A1(n5), .A2(n11), .ZN(B[11]) );
  CKND2D0BWP U21 ( .A1(A[3]), .A2(A[0]), .ZN(n5) );
  NR2D0BWP U22 ( .A1(n6), .A2(n11), .ZN(B[10]) );
  IND3D0BWP U23 ( .A1(A[4]), .B1(n3), .B2(A[1]), .ZN(n11) );
  CKND2D0BWP U24 ( .A1(A[3]), .A2(n2), .ZN(n6) );
  NR2D0BWP U25 ( .A1(n4), .A2(n9), .ZN(B[0]) );
  CKND2D0BWP U26 ( .A1(n2), .A2(n1), .ZN(n9) );
  OR3D0BWP U27 ( .A1(n12), .A2(A[1]), .A3(A[4]), .Z(n4) );
  NR2D0BWP U28 ( .A1(n3), .A2(A[4]), .ZN(n12) );
endmodule


module CVP14_DW01_add_1 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n2, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38;

  INVD1BWP U2 ( .I(n21), .ZN(n6) );
  INVD1BWP U3 ( .I(n29), .ZN(n7) );
  INVD1BWP U4 ( .I(n36), .ZN(n8) );
  INVD1BWP U5 ( .I(n38), .ZN(n9) );
  AN2XD1BWP U6 ( .A1(n2), .A2(n38), .Z(SUM[10]) );
  OR2XD1BWP U7 ( .A1(B[10]), .A2(A[10]), .Z(n2) );
  XOR2D1BWP U8 ( .A1(B[19]), .A2(n10), .Z(SUM[19]) );
  INVD1BWP U9 ( .I(B[18]), .ZN(n5) );
  CKBD1BWP U10 ( .I(A[8]), .Z(SUM[8]) );
  CKBD1BWP U11 ( .I(A[9]), .Z(SUM[9]) );
  MOAI22D0BWP U12 ( .A1(n11), .A2(n5), .B1(n12), .B2(A[18]), .ZN(n10) );
  NR2D0BWP U13 ( .A1(A[18]), .A2(n12), .ZN(n11) );
  XOR3D0BWP U14 ( .A1(B[18]), .A2(A[18]), .A3(n12), .Z(SUM[18]) );
  AO22D0BWP U15 ( .A1(n13), .A2(A[17]), .B1(n14), .B2(B[17]), .Z(n12) );
  OR2D0BWP U16 ( .A1(A[17]), .A2(n13), .Z(n14) );
  XOR3D0BWP U17 ( .A1(B[17]), .A2(A[17]), .A3(n13), .Z(SUM[17]) );
  OAI21D0BWP U18 ( .A1(n15), .A2(n16), .B(n17), .ZN(n13) );
  CKXOR2D0BWP U19 ( .A1(n16), .A2(n18), .Z(SUM[16]) );
  IND2D0BWP U20 ( .A1(n15), .B1(n17), .ZN(n18) );
  CKND2D0BWP U21 ( .A1(B[16]), .A2(A[16]), .ZN(n17) );
  NR2D0BWP U22 ( .A1(B[16]), .A2(A[16]), .ZN(n15) );
  AOI21D0BWP U23 ( .A1(n6), .A2(n19), .B(n20), .ZN(n16) );
  CKXOR2D0BWP U24 ( .A1(n22), .A2(n19), .Z(SUM[15]) );
  OAI21D0BWP U25 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  NR2D0BWP U26 ( .A1(n20), .A2(n21), .ZN(n22) );
  NR2D0BWP U27 ( .A1(B[15]), .A2(A[15]), .ZN(n21) );
  AN2D0BWP U28 ( .A1(B[15]), .A2(A[15]), .Z(n20) );
  CKXOR2D0BWP U29 ( .A1(n24), .A2(n26), .Z(SUM[14]) );
  IND2D0BWP U30 ( .A1(n23), .B1(n25), .ZN(n26) );
  CKND2D0BWP U31 ( .A1(B[14]), .A2(A[14]), .ZN(n25) );
  NR2D0BWP U32 ( .A1(B[14]), .A2(A[14]), .ZN(n23) );
  AOI21D0BWP U33 ( .A1(n7), .A2(n27), .B(n28), .ZN(n24) );
  CKXOR2D0BWP U34 ( .A1(n30), .A2(n27), .Z(SUM[13]) );
  OAI21D0BWP U35 ( .A1(n31), .A2(n32), .B(n33), .ZN(n27) );
  NR2D0BWP U36 ( .A1(n28), .A2(n29), .ZN(n30) );
  NR2D0BWP U37 ( .A1(B[13]), .A2(A[13]), .ZN(n29) );
  AN2D0BWP U38 ( .A1(B[13]), .A2(A[13]), .Z(n28) );
  CKXOR2D0BWP U39 ( .A1(n32), .A2(n34), .Z(SUM[12]) );
  IND2D0BWP U40 ( .A1(n31), .B1(n33), .ZN(n34) );
  CKND2D0BWP U41 ( .A1(B[12]), .A2(A[12]), .ZN(n33) );
  NR2D0BWP U42 ( .A1(B[12]), .A2(A[12]), .ZN(n31) );
  AOI21D0BWP U43 ( .A1(n8), .A2(n9), .B(n35), .ZN(n32) );
  CKXOR2D0BWP U44 ( .A1(n37), .A2(n9), .Z(SUM[11]) );
  NR2D0BWP U45 ( .A1(n35), .A2(n36), .ZN(n37) );
  NR2D0BWP U46 ( .A1(B[11]), .A2(A[11]), .ZN(n36) );
  AN2D0BWP U47 ( .A1(B[11]), .A2(A[11]), .Z(n35) );
  CKND2D0BWP U48 ( .A1(B[10]), .A2(A[10]), .ZN(n38) );
endmodule


module CVP14_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [10:0] A;
  input [10:0] B;
  output [21:0] PRODUCT;
  input TC;
  wire   \*Logic0* , \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] ,
         \ab[10][5] , \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] ,
         \ab[10][0] , \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] ,
         \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] ,
         \ab[9][1] , \ab[9][0] , \ab[8][10] , \ab[8][9] , \ab[8][8] ,
         \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] , \ab[8][3] ,
         \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][10] , \ab[7][9] ,
         \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] , \ab[7][4] ,
         \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] , \ab[6][10] ,
         \ab[6][9] , \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] ,
         \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] ,
         \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] ,
         \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] ,
         \ab[5][0] , \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] ,
         \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] ,
         \ab[4][1] , \ab[4][0] , \ab[3][10] , \ab[3][9] , \ab[3][8] ,
         \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][10] , \ab[2][9] ,
         \ab[2][8] , \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] ,
         \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] , \ab[1][10] ,
         \ab[1][9] , \ab[1][8] , \ab[1][7] , \ab[1][6] , \ab[1][5] ,
         \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[0][10] ,
         \ab[0][9] , \ab[0][8] , \ab[0][7] , \ab[0][6] , \ab[0][5] ,
         \ab[0][4] , \ab[0][3] , \ab[0][2] , \CARRYB[10][9] , \CARRYB[10][8] ,
         \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] , \CARRYB[10][4] ,
         \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] , \CARRYB[10][0] ,
         \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] ,
         \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] ,
         \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][9] , \CARRYB[8][8] ,
         \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] , \CARRYB[8][4] ,
         \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] , \CARRYB[8][0] ,
         \CARRYB[7][9] , \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] ,
         \CARRYB[7][5] , \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] ,
         \CARRYB[7][1] , \CARRYB[7][0] , \CARRYB[6][9] , \CARRYB[6][8] ,
         \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] ,
         \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] ,
         \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] ,
         \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] ,
         \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][9] , \CARRYB[4][8] ,
         \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] , \CARRYB[4][4] ,
         \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] , \CARRYB[4][0] ,
         \CARRYB[3][9] , \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] ,
         \CARRYB[3][5] , \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] ,
         \CARRYB[3][1] , \CARRYB[3][0] , \CARRYB[2][9] , \CARRYB[2][8] ,
         \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] ,
         \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] ,
         \CARRYB[1][9] , \CARRYB[1][8] , \CARRYB[1][7] , \CARRYB[1][6] ,
         \CARRYB[1][5] , \CARRYB[1][4] , \CARRYB[1][3] , \CARRYB[1][2] ,
         \CARRYB[1][1] , \CARRYB[1][0] , \SUMB[10][9] , \SUMB[10][8] ,
         \SUMB[10][7] , \SUMB[10][6] , \SUMB[10][5] , \SUMB[10][4] ,
         \SUMB[10][3] , \SUMB[10][2] , \SUMB[10][1] , \SUMB[10][0] ,
         \SUMB[9][9] , \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] ,
         \SUMB[9][4] , \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][9] ,
         \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] , \SUMB[8][4] ,
         \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][9] , \SUMB[7][8] ,
         \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] ,
         \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] ,
         \SUMB[6][6] , \SUMB[6][5] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] ,
         \SUMB[6][1] , \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][9] ,
         \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] , \SUMB[3][4] ,
         \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][9] , \SUMB[2][8] ,
         \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] ,
         \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] ,
         \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] ,
         \SUMB[1][1] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] ,
         \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[7] , \A1[6] , \A1[5] ,
         \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] , \A2[18] , \A2[17] ,
         \A2[16] , \A2[15] , \A2[14] , \A2[13] , \A2[12] , \A2[11] , \A2[10] ,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;
  assign \ab[10][9]  = B[9];
  assign \ab[10][8]  = B[8];
  assign \ab[10][7]  = B[7];
  assign \ab[10][6]  = B[6];
  assign \ab[10][5]  = B[5];
  assign \ab[10][4]  = B[4];
  assign \ab[10][3]  = B[3];
  assign \ab[10][2]  = B[2];
  assign \ab[10][1]  = B[1];
  assign \ab[10][0]  = B[0];
  assign \ab[9][10]  = A[9];
  assign \ab[8][10]  = A[8];
  assign \ab[7][10]  = A[7];
  assign \ab[6][10]  = A[6];
  assign \ab[5][10]  = A[5];
  assign \ab[4][10]  = A[4];
  assign \ab[3][10]  = A[3];
  assign \ab[2][10]  = A[2];
  assign \ab[1][10]  = A[1];
  assign \ab[0][10]  = A[0];

  CVP14_DW01_add_1 FS_1 ( .A({\*Logic0* , n19, \A1[17] , \A1[16] , \A1[15] , 
        \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , 
        \SUMB[10][0] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , 
        \A1[1] , \A1[0] }), .B({\CARRYB[10][9] , \A2[18] , \A2[17] , \A2[16] , 
        \A2[15] , \A2[14] , \A2[13] , \A2[12] , \A2[11] , \A2[10] , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* }), .CI(\*Logic0* ), .SUM({
        PRODUCT[21:10], SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7}) );
  FA1D0BWP S3_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\ab[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA1D0BWP S3_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\ab[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA1D0BWP S3_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\ab[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA1D0BWP S3_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\ab[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA1D0BWP S3_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\ab[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA1D0BWP S3_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\ab[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA1D0BWP S3_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\ab[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA1D0BWP S2_2_8 ( .A(\ab[2][8] ), .B(\CARRYB[1][8] ), .CI(\SUMB[1][9] ), 
        .CO(\CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FA1D0BWP S3_2_9 ( .A(\ab[2][9] ), .B(\CARRYB[1][9] ), .CI(\ab[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FA1D0BWP S5_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\ab[9][10] ), .CO(
        \CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA1D0BWP S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), 
        .CO(\CARRYB[8][0] ), .S(\A1[6] ) );
  FA1D0BWP S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), 
        .CO(\CARRYB[9][0] ), .S(\A1[7] ) );
  FA1D0BWP S4_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\SUMB[10][0] ) );
  FA1D0BWP S4_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA1D0BWP S4_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA1D0BWP S4_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA1D0BWP S4_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA1D0BWP S4_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA1D0BWP S4_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA1D0BWP S4_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA1D0BWP S4_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA1D0BWP S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), 
        .CO(\CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA1D0BWP S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), 
        .CO(\CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA1D0BWP S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), 
        .CO(\CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA1D0BWP S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), 
        .CO(\CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA1D0BWP S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), 
        .CO(\CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA1D0BWP S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), 
        .CO(\CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA1D0BWP S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), 
        .CO(\CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA1D0BWP S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), 
        .CO(\CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA1D0BWP S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), 
        .CO(\CARRYB[5][0] ), .S(\A1[3] ) );
  FA1D0BWP S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), 
        .CO(\CARRYB[6][0] ), .S(\A1[4] ) );
  FA1D0BWP S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), 
        .CO(\CARRYB[7][0] ), .S(\A1[5] ) );
  FA1D0BWP S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), 
        .CO(\CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA1D0BWP S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), 
        .CO(\CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA1D0BWP S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), 
        .CO(\CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA1D0BWP S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), 
        .CO(\CARRYB[2][0] ), .S(\A1[0] ) );
  FA1D0BWP S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), 
        .CO(\CARRYB[3][0] ), .S(\A1[1] ) );
  FA1D0BWP S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), 
        .CO(\CARRYB[4][0] ), .S(\A1[2] ) );
  FA1D0BWP S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), 
        .CO(\CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA1D0BWP S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), 
        .CO(\CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA1D0BWP S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), 
        .CO(\CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA1D0BWP S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), 
        .CO(\CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA1D0BWP S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), 
        .CO(\CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA1D0BWP S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), 
        .CO(\CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA1D0BWP S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), 
        .CO(\CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA1D0BWP S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), 
        .CO(\CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA1D0BWP S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), 
        .CO(\CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA1D0BWP S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), 
        .CO(\CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA1D0BWP S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), 
        .CO(\CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA1D0BWP S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), 
        .CO(\CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA1D0BWP S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), 
        .CO(\CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA1D0BWP S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), 
        .CO(\CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA1D0BWP S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), 
        .CO(\CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA1D0BWP S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), 
        .CO(\CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA1D0BWP S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), 
        .CO(\CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA1D0BWP S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), 
        .CO(\CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA1D0BWP S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), 
        .CO(\CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA1D0BWP S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), 
        .CO(\CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA1D0BWP S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), 
        .CO(\CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA1D0BWP S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), 
        .CO(\CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA1D0BWP S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), 
        .CO(\CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA1D0BWP S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), 
        .CO(\CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA1D0BWP S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), 
        .CO(\CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA1D0BWP S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), 
        .CO(\CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA1D0BWP S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), 
        .CO(\CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA1D0BWP S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), 
        .CO(\CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA1D0BWP S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), 
        .CO(\CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA1D0BWP S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), 
        .CO(\CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA1D0BWP S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), 
        .CO(\CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA1D0BWP S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), 
        .CO(\CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA1D0BWP S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), 
        .CO(\CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA1D0BWP S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), 
        .CO(\CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA1D0BWP S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), 
        .CO(\CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA1D0BWP S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), 
        .CO(\CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA1D0BWP S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), 
        .CO(\CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA1D0BWP S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), 
        .CO(\CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA1D0BWP S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), 
        .CO(\CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA1D0BWP S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), 
        .CO(\CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA1D0BWP S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), 
        .CO(\CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA1D0BWP S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), 
        .CO(\CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA1D0BWP S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), 
        .CO(\CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA1D0BWP S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), 
        .CO(\CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA1D0BWP S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), 
        .CO(\CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA1D0BWP S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), 
        .CO(\CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FA1D0BWP S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), 
        .CO(\CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FA1D0BWP S2_2_3 ( .A(\ab[2][3] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), 
        .CO(\CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FA1D0BWP S2_2_4 ( .A(\ab[2][4] ), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), 
        .CO(\CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FA1D0BWP S2_2_5 ( .A(\ab[2][5] ), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), 
        .CO(\CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FA1D0BWP S2_2_6 ( .A(\ab[2][6] ), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), 
        .CO(\CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FA1D0BWP S2_2_7 ( .A(\ab[2][7] ), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), 
        .CO(\CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  INVD1BWP U2 ( .I(\ab[0][7] ), .ZN(n13) );
  INVD1BWP U3 ( .I(\ab[0][6] ), .ZN(n11) );
  INVD1BWP U4 ( .I(\ab[0][5] ), .ZN(n9) );
  INVD1BWP U5 ( .I(\ab[0][4] ), .ZN(n7) );
  INVD1BWP U6 ( .I(\ab[0][3] ), .ZN(n5) );
  INVD1BWP U7 ( .I(\ab[0][2] ), .ZN(n3) );
  INVD1BWP U8 ( .I(\ab[0][9] ), .ZN(n17) );
  INVD1BWP U9 ( .I(\ab[0][8] ), .ZN(n15) );
  INVD1BWP U10 ( .I(\ab[1][1] ), .ZN(n2) );
  INVD1BWP U11 ( .I(\ab[1][7] ), .ZN(n14) );
  INVD1BWP U12 ( .I(\ab[1][6] ), .ZN(n12) );
  INVD1BWP U13 ( .I(\ab[1][5] ), .ZN(n10) );
  INVD1BWP U14 ( .I(\ab[1][4] ), .ZN(n8) );
  INVD1BWP U15 ( .I(\ab[1][3] ), .ZN(n6) );
  INVD1BWP U16 ( .I(\ab[1][2] ), .ZN(n4) );
  INVD1BWP U17 ( .I(\ab[1][9] ), .ZN(n18) );
  INVD1BWP U18 ( .I(\ab[1][8] ), .ZN(n16) );
  CKXOR2D0BWP U19 ( .A1(\ab[1][1] ), .A2(\ab[0][2] ), .Z(\SUMB[1][1] ) );
  NR2XD0BWP U20 ( .A1(n14), .A2(n15), .ZN(\CARRYB[1][7] ) );
  CKXOR2D0BWP U21 ( .A1(\ab[1][8] ), .A2(\ab[0][9] ), .Z(\SUMB[1][8] ) );
  NR2XD0BWP U22 ( .A1(n12), .A2(n13), .ZN(\CARRYB[1][6] ) );
  CKXOR2D0BWP U23 ( .A1(\ab[1][7] ), .A2(\ab[0][8] ), .Z(\SUMB[1][7] ) );
  NR2XD0BWP U24 ( .A1(n10), .A2(n11), .ZN(\CARRYB[1][5] ) );
  CKXOR2D0BWP U25 ( .A1(\ab[1][6] ), .A2(\ab[0][7] ), .Z(\SUMB[1][6] ) );
  NR2XD0BWP U26 ( .A1(n8), .A2(n9), .ZN(\CARRYB[1][4] ) );
  CKXOR2D0BWP U27 ( .A1(\ab[1][5] ), .A2(\ab[0][6] ), .Z(\SUMB[1][5] ) );
  NR2XD0BWP U28 ( .A1(n6), .A2(n7), .ZN(\CARRYB[1][3] ) );
  CKXOR2D0BWP U29 ( .A1(\ab[1][4] ), .A2(\ab[0][5] ), .Z(\SUMB[1][4] ) );
  NR2XD0BWP U30 ( .A1(n4), .A2(n5), .ZN(\CARRYB[1][2] ) );
  CKXOR2D0BWP U31 ( .A1(\ab[1][3] ), .A2(\ab[0][4] ), .Z(\SUMB[1][3] ) );
  NR2XD0BWP U32 ( .A1(n2), .A2(n3), .ZN(\CARRYB[1][1] ) );
  CKXOR2D0BWP U33 ( .A1(\ab[1][2] ), .A2(\ab[0][3] ), .Z(\SUMB[1][2] ) );
  XOR2D1BWP U34 ( .A1(\SUMB[10][9] ), .A2(\CARRYB[10][8] ), .Z(\A1[17] ) );
  XOR2D1BWP U35 ( .A1(\SUMB[10][3] ), .A2(\CARRYB[10][2] ), .Z(\A1[11] ) );
  XOR2D1BWP U36 ( .A1(\SUMB[10][5] ), .A2(\CARRYB[10][4] ), .Z(\A1[13] ) );
  XOR2D1BWP U37 ( .A1(\SUMB[10][7] ), .A2(\CARRYB[10][6] ), .Z(\A1[15] ) );
  XOR2D1BWP U38 ( .A1(\SUMB[10][4] ), .A2(\CARRYB[10][3] ), .Z(\A1[12] ) );
  XOR2D1BWP U39 ( .A1(\SUMB[10][6] ), .A2(\CARRYB[10][5] ), .Z(\A1[14] ) );
  XOR2D1BWP U40 ( .A1(\SUMB[10][8] ), .A2(\CARRYB[10][7] ), .Z(\A1[16] ) );
  XOR2D1BWP U41 ( .A1(\SUMB[10][2] ), .A2(\CARRYB[10][1] ), .Z(\A1[10] ) );
  XOR2D1BWP U42 ( .A1(\SUMB[10][1] ), .A2(\CARRYB[10][0] ), .Z(\A1[9] ) );
  AN2XD1BWP U43 ( .A1(\CARRYB[10][8] ), .A2(\SUMB[10][9] ), .Z(\A2[18] ) );
  INVD1BWP U44 ( .I(\CARRYB[10][9] ), .ZN(n19) );
  AN2XD1BWP U45 ( .A1(\CARRYB[10][7] ), .A2(\SUMB[10][8] ), .Z(\A2[17] ) );
  AN2XD1BWP U46 ( .A1(\CARRYB[10][1] ), .A2(\SUMB[10][2] ), .Z(\A2[11] ) );
  AN2XD1BWP U47 ( .A1(\CARRYB[10][3] ), .A2(\SUMB[10][4] ), .Z(\A2[13] ) );
  AN2XD1BWP U48 ( .A1(\CARRYB[10][5] ), .A2(\SUMB[10][6] ), .Z(\A2[15] ) );
  AN2XD1BWP U49 ( .A1(\CARRYB[10][2] ), .A2(\SUMB[10][3] ), .Z(\A2[12] ) );
  AN2XD1BWP U50 ( .A1(\CARRYB[10][4] ), .A2(\SUMB[10][5] ), .Z(\A2[14] ) );
  AN2XD1BWP U51 ( .A1(\CARRYB[10][6] ), .A2(\SUMB[10][7] ), .Z(\A2[16] ) );
  AN2XD1BWP U52 ( .A1(\CARRYB[10][0] ), .A2(\SUMB[10][1] ), .Z(\A2[10] ) );
  NR2XD0BWP U53 ( .A1(n18), .A2(n39), .ZN(\CARRYB[1][9] ) );
  NR2XD0BWP U54 ( .A1(n16), .A2(n17), .ZN(\CARRYB[1][8] ) );
  CKXOR2D0BWP U55 ( .A1(\ab[1][9] ), .A2(\ab[0][10] ), .Z(\SUMB[1][9] ) );
  INVD1BWP U56 ( .I(\ab[0][10] ), .ZN(n39) );
  INVD1BWP U57 ( .I(\ab[10][7] ), .ZN(n22) );
  INVD1BWP U58 ( .I(\ab[10][3] ), .ZN(n26) );
  INVD1BWP U59 ( .I(\ab[10][4] ), .ZN(n25) );
  INVD1BWP U60 ( .I(\ab[10][6] ), .ZN(n23) );
  INVD1BWP U61 ( .I(\ab[10][5] ), .ZN(n24) );
  INVD1BWP U62 ( .I(\ab[3][10] ), .ZN(n31) );
  INVD1BWP U63 ( .I(\ab[5][10] ), .ZN(n34) );
  INVD1BWP U64 ( .I(\ab[4][10] ), .ZN(n30) );
  INVD1BWP U65 ( .I(\ab[6][10] ), .ZN(n35) );
  INVD1BWP U66 ( .I(\ab[10][2] ), .ZN(n27) );
  INVD1BWP U67 ( .I(\ab[2][10] ), .ZN(n32) );
  INVD1BWP U68 ( .I(\ab[7][10] ), .ZN(n36) );
  INVD1BWP U69 ( .I(\ab[10][1] ), .ZN(n28) );
  INVD1BWP U70 ( .I(\ab[10][0] ), .ZN(n29) );
  INVD1BWP U71 ( .I(\ab[1][10] ), .ZN(n33) );
  INVD1BWP U72 ( .I(\ab[8][10] ), .ZN(n37) );
  INVD1BWP U73 ( .I(\ab[9][10] ), .ZN(n38) );
  INVD1BWP U74 ( .I(\ab[10][8] ), .ZN(n21) );
  INVD1BWP U75 ( .I(\ab[10][9] ), .ZN(n20) );
  TIELBWP U76 ( .ZN(\*Logic0* ) );
  NR2D0BWP U77 ( .A1(n38), .A2(n20), .ZN(\ab[9][9] ) );
  NR2D0BWP U78 ( .A1(n38), .A2(n21), .ZN(\ab[9][8] ) );
  NR2D0BWP U79 ( .A1(n38), .A2(n22), .ZN(\ab[9][7] ) );
  NR2D0BWP U80 ( .A1(n38), .A2(n23), .ZN(\ab[9][6] ) );
  NR2D0BWP U81 ( .A1(n38), .A2(n24), .ZN(\ab[9][5] ) );
  NR2D0BWP U82 ( .A1(n38), .A2(n25), .ZN(\ab[9][4] ) );
  NR2D0BWP U83 ( .A1(n38), .A2(n26), .ZN(\ab[9][3] ) );
  NR2D0BWP U84 ( .A1(n38), .A2(n27), .ZN(\ab[9][2] ) );
  NR2D0BWP U85 ( .A1(n38), .A2(n28), .ZN(\ab[9][1] ) );
  NR2D0BWP U86 ( .A1(n38), .A2(n29), .ZN(\ab[9][0] ) );
  NR2D0BWP U87 ( .A1(n20), .A2(n37), .ZN(\ab[8][9] ) );
  NR2D0BWP U88 ( .A1(n21), .A2(n37), .ZN(\ab[8][8] ) );
  NR2D0BWP U89 ( .A1(n22), .A2(n37), .ZN(\ab[8][7] ) );
  NR2D0BWP U90 ( .A1(n23), .A2(n37), .ZN(\ab[8][6] ) );
  NR2D0BWP U91 ( .A1(n24), .A2(n37), .ZN(\ab[8][5] ) );
  NR2D0BWP U92 ( .A1(n25), .A2(n37), .ZN(\ab[8][4] ) );
  NR2D0BWP U93 ( .A1(n26), .A2(n37), .ZN(\ab[8][3] ) );
  NR2D0BWP U94 ( .A1(n27), .A2(n37), .ZN(\ab[8][2] ) );
  NR2D0BWP U95 ( .A1(n28), .A2(n37), .ZN(\ab[8][1] ) );
  NR2D0BWP U96 ( .A1(n29), .A2(n37), .ZN(\ab[8][0] ) );
  NR2D0BWP U97 ( .A1(n20), .A2(n36), .ZN(\ab[7][9] ) );
  NR2D0BWP U98 ( .A1(n21), .A2(n36), .ZN(\ab[7][8] ) );
  NR2D0BWP U99 ( .A1(n22), .A2(n36), .ZN(\ab[7][7] ) );
  NR2D0BWP U100 ( .A1(n23), .A2(n36), .ZN(\ab[7][6] ) );
  NR2D0BWP U101 ( .A1(n24), .A2(n36), .ZN(\ab[7][5] ) );
  NR2D0BWP U102 ( .A1(n25), .A2(n36), .ZN(\ab[7][4] ) );
  NR2D0BWP U103 ( .A1(n26), .A2(n36), .ZN(\ab[7][3] ) );
  NR2D0BWP U104 ( .A1(n27), .A2(n36), .ZN(\ab[7][2] ) );
  NR2D0BWP U105 ( .A1(n28), .A2(n36), .ZN(\ab[7][1] ) );
  NR2D0BWP U106 ( .A1(n29), .A2(n36), .ZN(\ab[7][0] ) );
  NR2D0BWP U107 ( .A1(n20), .A2(n35), .ZN(\ab[6][9] ) );
  NR2D0BWP U108 ( .A1(n21), .A2(n35), .ZN(\ab[6][8] ) );
  NR2D0BWP U109 ( .A1(n22), .A2(n35), .ZN(\ab[6][7] ) );
  NR2D0BWP U110 ( .A1(n23), .A2(n35), .ZN(\ab[6][6] ) );
  NR2D0BWP U111 ( .A1(n24), .A2(n35), .ZN(\ab[6][5] ) );
  NR2D0BWP U112 ( .A1(n25), .A2(n35), .ZN(\ab[6][4] ) );
  NR2D0BWP U113 ( .A1(n26), .A2(n35), .ZN(\ab[6][3] ) );
  NR2D0BWP U114 ( .A1(n27), .A2(n35), .ZN(\ab[6][2] ) );
  NR2D0BWP U115 ( .A1(n28), .A2(n35), .ZN(\ab[6][1] ) );
  NR2D0BWP U116 ( .A1(n29), .A2(n35), .ZN(\ab[6][0] ) );
  NR2D0BWP U117 ( .A1(n20), .A2(n34), .ZN(\ab[5][9] ) );
  NR2D0BWP U118 ( .A1(n21), .A2(n34), .ZN(\ab[5][8] ) );
  NR2D0BWP U119 ( .A1(n22), .A2(n34), .ZN(\ab[5][7] ) );
  NR2D0BWP U120 ( .A1(n23), .A2(n34), .ZN(\ab[5][6] ) );
  NR2D0BWP U121 ( .A1(n24), .A2(n34), .ZN(\ab[5][5] ) );
  NR2D0BWP U122 ( .A1(n25), .A2(n34), .ZN(\ab[5][4] ) );
  NR2D0BWP U123 ( .A1(n26), .A2(n34), .ZN(\ab[5][3] ) );
  NR2D0BWP U124 ( .A1(n27), .A2(n34), .ZN(\ab[5][2] ) );
  NR2D0BWP U125 ( .A1(n28), .A2(n34), .ZN(\ab[5][1] ) );
  NR2D0BWP U126 ( .A1(n29), .A2(n34), .ZN(\ab[5][0] ) );
  NR2D0BWP U127 ( .A1(n20), .A2(n30), .ZN(\ab[4][9] ) );
  NR2D0BWP U128 ( .A1(n21), .A2(n30), .ZN(\ab[4][8] ) );
  NR2D0BWP U129 ( .A1(n22), .A2(n30), .ZN(\ab[4][7] ) );
  NR2D0BWP U130 ( .A1(n23), .A2(n30), .ZN(\ab[4][6] ) );
  NR2D0BWP U131 ( .A1(n24), .A2(n30), .ZN(\ab[4][5] ) );
  NR2D0BWP U132 ( .A1(n25), .A2(n30), .ZN(\ab[4][4] ) );
  NR2D0BWP U133 ( .A1(n26), .A2(n30), .ZN(\ab[4][3] ) );
  NR2D0BWP U134 ( .A1(n27), .A2(n30), .ZN(\ab[4][2] ) );
  NR2D0BWP U135 ( .A1(n28), .A2(n30), .ZN(\ab[4][1] ) );
  NR2D0BWP U136 ( .A1(n29), .A2(n30), .ZN(\ab[4][0] ) );
  NR2D0BWP U137 ( .A1(n20), .A2(n31), .ZN(\ab[3][9] ) );
  NR2D0BWP U138 ( .A1(n21), .A2(n31), .ZN(\ab[3][8] ) );
  NR2D0BWP U139 ( .A1(n22), .A2(n31), .ZN(\ab[3][7] ) );
  NR2D0BWP U140 ( .A1(n23), .A2(n31), .ZN(\ab[3][6] ) );
  NR2D0BWP U141 ( .A1(n24), .A2(n31), .ZN(\ab[3][5] ) );
  NR2D0BWP U142 ( .A1(n25), .A2(n31), .ZN(\ab[3][4] ) );
  NR2D0BWP U143 ( .A1(n26), .A2(n31), .ZN(\ab[3][3] ) );
  NR2D0BWP U144 ( .A1(n27), .A2(n31), .ZN(\ab[3][2] ) );
  NR2D0BWP U145 ( .A1(n28), .A2(n31), .ZN(\ab[3][1] ) );
  NR2D0BWP U146 ( .A1(n29), .A2(n31), .ZN(\ab[3][0] ) );
  NR2D0BWP U147 ( .A1(n20), .A2(n32), .ZN(\ab[2][9] ) );
  NR2D0BWP U148 ( .A1(n21), .A2(n32), .ZN(\ab[2][8] ) );
  NR2D0BWP U149 ( .A1(n22), .A2(n32), .ZN(\ab[2][7] ) );
  NR2D0BWP U150 ( .A1(n23), .A2(n32), .ZN(\ab[2][6] ) );
  NR2D0BWP U151 ( .A1(n24), .A2(n32), .ZN(\ab[2][5] ) );
  NR2D0BWP U152 ( .A1(n25), .A2(n32), .ZN(\ab[2][4] ) );
  NR2D0BWP U153 ( .A1(n26), .A2(n32), .ZN(\ab[2][3] ) );
  NR2D0BWP U154 ( .A1(n27), .A2(n32), .ZN(\ab[2][2] ) );
  NR2D0BWP U155 ( .A1(n28), .A2(n32), .ZN(\ab[2][1] ) );
  NR2D0BWP U156 ( .A1(n29), .A2(n32), .ZN(\ab[2][0] ) );
  NR2D0BWP U157 ( .A1(n20), .A2(n33), .ZN(\ab[1][9] ) );
  NR2D0BWP U158 ( .A1(n21), .A2(n33), .ZN(\ab[1][8] ) );
  NR2D0BWP U159 ( .A1(n22), .A2(n33), .ZN(\ab[1][7] ) );
  NR2D0BWP U160 ( .A1(n23), .A2(n33), .ZN(\ab[1][6] ) );
  NR2D0BWP U161 ( .A1(n24), .A2(n33), .ZN(\ab[1][5] ) );
  NR2D0BWP U162 ( .A1(n25), .A2(n33), .ZN(\ab[1][4] ) );
  NR2D0BWP U163 ( .A1(n26), .A2(n33), .ZN(\ab[1][3] ) );
  NR2D0BWP U164 ( .A1(n27), .A2(n33), .ZN(\ab[1][2] ) );
  NR2D0BWP U165 ( .A1(n20), .A2(n39), .ZN(\ab[0][9] ) );
  NR2D0BWP U166 ( .A1(n21), .A2(n39), .ZN(\ab[0][8] ) );
  NR2D0BWP U167 ( .A1(n22), .A2(n39), .ZN(\ab[0][7] ) );
  NR2D0BWP U168 ( .A1(n23), .A2(n39), .ZN(\ab[0][6] ) );
  NR2D0BWP U169 ( .A1(n24), .A2(n39), .ZN(\ab[0][5] ) );
  NR2D0BWP U170 ( .A1(n25), .A2(n39), .ZN(\ab[0][4] ) );
  NR2D0BWP U171 ( .A1(n26), .A2(n39), .ZN(\ab[0][3] ) );
  NR2D0BWP U172 ( .A1(n27), .A2(n39), .ZN(\ab[0][2] ) );
  AN3D0BWP U173 ( .A1(\ab[1][1] ), .A2(\ab[10][0] ), .A3(\ab[0][10] ), .Z(
        \CARRYB[1][0] ) );
  NR2D0BWP U174 ( .A1(n33), .A2(n28), .ZN(\ab[1][1] ) );
endmodule


module CVP14 ( Addr, RD, WR, V, dataOut, Reset, Clk1, Clk2, DataIn );
  output [15:0] Addr;
  output [15:0] dataOut;
  input [15:0] DataIn;
  input Reset, Clk1, Clk2;
  output RD, WR, V;
  wire   N137, N138, N139, N140, overflow, N207, N208, N209, N210, N211, N212,
         N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N253,
         N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264,
         N265, N266, N267, N317, N318, N319, N320, N321, N322, N323, N324,
         N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335,
         N336, N337, N338, N339, N340, N341, N342, N343, N344, N345, N346,
         N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, N357,
         N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368,
         N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N401,
         N402, N403, N404, N405, N406, N407, N408, N409, N410, N411, N412,
         N413, N414, N415, N416, N417, N418, N419, N420, N421, N422, N423,
         N424, N425, N426, N427, N428, N429, N430, N431, N432, N433, N434,
         N435, N436, N437, N438, N439, N440, N441, N442, N443, N444, N445,
         N446, N447, N448, N449, N450, N451, N452, N453, N454, N455, N456,
         N457, N458, N459, N460, N461, N462, N463, N464, N465, N466, N467,
         N468, N469, N470, N471, N472, N473, N474, N475, N476, N477, N478,
         N479, N480, N481, N482, N483, N484, N485, N486, N487, N488, N489,
         N490, N491, N492, N493, N494, N495, N496, N497, N498, N499, N500,
         N501, N502, N503, N504, N505, N506, N507, N508, N509, N510, N511,
         N512, N513, N514, N515, N516, N517, N518, N519, N520, N521, N522,
         N523, N524, N525, N526, N527, N528, N529, N530, N531, N532, N533,
         N534, N535, N536, N537, N538, N539, N540, N541, N542, N543, N544,
         N545, N546, N547, N548, N549, N550, N551, N552, N553, N554, N555,
         N556, N557, N558, N559, N560, N561, N562, N563, N564, N565, N566,
         N567, N568, N569, N570, N571, N572, N1094, N1095, N1096, N1097, N1098,
         N1099, N1100, N1101, N1102, N1103, N1104, N1105, N1106, N1107, N1108,
         N1163, N1164, N1165, N1166, N1167, N1168, N1169, N1173, N1174, N1175,
         N1176, N1177, N1178, N1179, N1180, N1181, N1182, N1183, N1184, N1185,
         N1186, N1187, N1188, N1189, N1190, N1191, N1192, N1193, N1194, N1195,
         N1196, N1197, N1198, N1254, N1255, N1256, N1257, N1258, N1259, N1260,
         N1261, N1262, N1263, N1264, N1265, N1266, N1280, N1282, N1283, N1284,
         N1285, N1286, N1287, N1288, N1289, N1290, N1291, N1292, N1293, N1294,
         N1295, N1296, N1297, N1298, N1299, N1300, N1301, N1302, N1303, N1304,
         N1305, N1306, N1307, N1407, N1408, N1409, N1410, N1411, N1412, N1413,
         N1414, N1415, N1416, N1417, N1418, N1419, N1457, N1466, N1487, N1488,
         N1489, N1490, N1491, N1492, N1493, N1494, N1495, N1496, N1497, N1498,
         N1499, N1500, N1512, N1513, N1514, N1519, N1520, N1521, N1522, N1523,
         N1524, N1527, N1528, N1529, N1530, N1531, N1532, N1533, N1534, N1535,
         N1536, N1537, N1545, N1546, N1547, N1548, N1549, N1550, N1551, N1552,
         N1553, N1554, N1555, N1556, N1557, N1558, N1561, N1562, N1563, N1564,
         N1565, N1600, N1601, N1602, N1610, N1660, N1681, N1682, N1683, N1684,
         N1685, N1686, N1687, N1688, N1689, N1690, N1691, N1747, N1748, N1749,
         N1750, N1751, N1752, N1753, N1754, N1755, N1756, N1757, N1758, N1759,
         N1760, N1761, N1762, N1772, N1773, N1774, N1775, N1776, N1777, N1778,
         N1779, N1780, N1781, N1782, N1783, N1784, N1785, N1786, N2626, N2627,
         N2628, N2629, N2630, N2631, N2632, N2633, N2634, N2635, N2636, N2637,
         N2638, N2639, N2640, N2641, N2642, N2643, N2644, N2645, N2646, N2647,
         N2648, N2649, N2650, N2651, N2652, N2653, N2654, N2655, N2656, N2657,
         N2658, N2659, N2660, N2661, N2662, N2663, N2664, N2665, N2666, N2667,
         N2668, N2669, N2670, N2671, N2672, N2673, N2674, N2675, N2676, N2677,
         N2678, N2679, N2680, N2681, N2682, N2683, N2684, N2685, N2686, N2687,
         N2688, N2689, N2690, N2691, N2692, N2693, N2694, N2695, N2696, N2697,
         N2698, N2699, N2700, N2701, N2702, N2703, N2704, N2705, N2706, N2707,
         N2708, N2709, N2710, N2711, N2712, N2713, N2714, N2715, N2716, N2717,
         N2718, N2719, N2720, N2721, N2722, N2723, N2724, N2725, N2726, N2727,
         N2728, N2729, N2730, N2731, N2732, N2733, N2734, N2735, N2736, N2737,
         N2738, N2739, N2740, N2741, N2742, N2743, N2744, N2745, N2746, N2747,
         N2748, N2749, N2750, N2751, N2752, N2753, N2754, N2755, N2756, N2757,
         N2758, N2759, N2760, N2761, N2762, N2763, N2764, N2765, N2766, N2767,
         N2768, N2769, N2770, N2771, N2772, N2773, N2774, N2775, N2776, N2777,
         N2778, N2779, N2780, N2781, N2782, N2783, N2784, N2785, N2786, N2787,
         N2788, N2789, N2790, N2791, N2792, N2793, N2794, N2795, N2796, N2797,
         N2798, N2799, N2800, N2801, N2802, N2803, N2804, N2805, N2806, N2807,
         N2808, N2809, N2810, N2811, N2812, N2813, N2814, N2815, N2816, N2817,
         N2818, N2819, N2820, N2821, N2822, N2823, N2824, N2825, N2826, N2827,
         N2828, N2829, N2830, N2831, N2832, N2833, N2834, N2835, N2836, N2837,
         N2838, N2839, N2840, N2841, N2842, N2843, N2844, N2845, N2846, N2847,
         N2848, N2849, N2850, N2851, N2852, N2853, N2854, N2855, N2856, N2857,
         N2858, N2859, N2860, N2861, N2862, N2863, N2864, N2865, N2866, N2867,
         N2868, N2869, N2870, N2871, N2872, N2873, N2874, N2875, N2876, N2877,
         N2878, N2879, N2880, N2881, N2882, N3432, N3433, N3434, N3435, N3436,
         N3753, N3754, N3755, N3756, N3757, N3758, N3759, N3760, N3761, N3762,
         N3763, N3764, N3765, N3766, N3767, N3768, N4028, N4029, N4030, N4031,
         N4032, N4033, N4034, N4035, N4036, N4037, N4038, N4039, N4040, N4041,
         N4042, N4043, N4044, N4047, N4048, N4049, N4050, N4051, N4052, N4053,
         N4054, N4055, N4056, N4057, N4058, N4059, N4060, N4061, N4062, N4063,
         N4064, N4065, N4066, N4067, N4068, N4069, N4070, N4071, N4072, N4073,
         N4074, N4075, N4076, N4077, N4078, N4079, N4080, N4081, N4082, N4083,
         N4084, N4085, N4086, N4087, N4088, N4089, N4090, N4091, N4092, N4093,
         N4094, N4095, N4096, N4097, N4098, N4099, N4100, N4101, N4102, N4103,
         N4104, N4105, N4106, N4107, N4108, N4109, N4110, N4111, N4112, N4113,
         N4114, N4115, N4116, N4117, N4118, N4119, N4120, N4121, N4123, N4124,
         N4125, N4126, N4127, N4128, N4129, N4130, N4131, N4132, N4133, N4134,
         N4135, N4136, N4137, N4138, N4139, N4140, N4141, N4142, N4143, N4144,
         N4145, N4146, N4147, N4148, N4149, N4150, N4151, N4152, N4153, N4154,
         N4155, N4156, N4157, N4158, N4159, N4160, N4161, N4162, N4163, N4164,
         N4165, N4166, N4167, N4168, N4169, N4170, N4171, N4172, N4173, N4174,
         N4175, N4176, N4177, N4178, N4179, N4180, N4181, N4182, N4183, N4184,
         N4185, N4186, N4187, N4188, N4189, N4190, N4191, N4192, N4193, N4194,
         N4195, N4196, N4197, N4198, N4199, N4200, N4201, N4202, N4203, N4204,
         N4205, N4206, N4207, N4208, N4209, N4210, N4211, N4212, N4213, N4214,
         N4215, N4216, N4217, N4218, N4219, N4220, N4221, N4223, N4224, N4225,
         N4226, N4227, N4228, N4229, N4230, N4231, N4232, N4233, N4234, N4235,
         N4236, N4237, N4238, N4239, N4240, N4241, N4242, N4243, N4244, N4245,
         N4246, N4247, N4248, N4249, N4250, N4251, N4252, N4253, N4254, N4255,
         N4256, N4257, N4258, N4259, N4260, N4261, N4262, N4263, N4264, N4265,
         N4266, N4267, N4268, N4269, N4270, N4271, N4272, N4273, N4274, N4275,
         N4276, N4277, N4278, N4279, N4280, N4281, N4282, N4283, N4284, N4285,
         N4286, N4287, N4288, N4289, N4290, N4291, N4292, N4293, N4294, N4295,
         N4296, N4297, N4298, N4299, N4300, N4301, N4302, N4303, N4304, N4305,
         N4306, N4307, N4308, N4309, N4310, N4311, N4312, N4313, N4314, N4315,
         N4316, N4317, N4318, N4319, N4320, N4321, N4322, N4323, N4324, N4325,
         N4326, N4327, N4328, N4329, N4330, N4331, N4332, N4333, N4334, N4335,
         N4336, N4337, N4338, N4339, N4340, N4341, N4342, N4343, N4344, N4345,
         N4346, N4347, N4348, N4349, N4350, N4351, N4352, N4353, N4354, N4355,
         N4356, N4357, N4358, N4359, N4360, N4361, N4362, N4363, N4364, N4366,
         \vrf/N296 , \vrf/N293 , \vrf/N290 , \vrf/N287 , \vrf/N284 ,
         \vrf/N281 , \vrf/N278 , \vrf/N275 , \vrf/N274 , \vrf/N273 ,
         \vrf/N272 , \vrf/N271 , \vrf/N270 , \vrf/N269 , \vrf/N268 ,
         \vrf/N267 , \vrf/N266 , \vrf/N265 , \vrf/N264 , \vrf/N263 ,
         \vrf/N262 , \vrf/N261 , \vrf/N260 , \vrf/N259 , \vrf/N258 ,
         \vrf/N257 , \vrf/N256 , \vrf/N255 , \vrf/N254 , \vrf/N253 ,
         \vrf/N252 , \vrf/N251 , \vrf/N250 , \vrf/N249 , \vrf/N248 ,
         \vrf/N247 , \vrf/N246 , \vrf/N245 , \vrf/N244 , \vrf/N243 ,
         \vrf/N242 , \vrf/N241 , \vrf/N240 , \vrf/N239 , \vrf/N238 ,
         \vrf/N237 , \vrf/N236 , \vrf/N235 , \vrf/N234 , \vrf/N233 ,
         \vrf/N232 , \vrf/N231 , \vrf/N230 , \vrf/N229 , \vrf/N228 ,
         \vrf/N227 , \vrf/N226 , \vrf/N225 , \vrf/N224 , \vrf/N223 ,
         \vrf/N222 , \vrf/N221 , \vrf/N220 , \vrf/N219 , \vrf/N218 ,
         \vrf/N217 , \vrf/N216 , \vrf/N215 , \vrf/N214 , \vrf/N213 ,
         \vrf/N212 , \vrf/N211 , \vrf/N210 , \vrf/N209 , \vrf/N208 ,
         \vrf/N207 , \vrf/N206 , \vrf/N205 , \vrf/N204 , \vrf/N203 ,
         \vrf/N202 , \vrf/N201 , \vrf/N200 , \vrf/N199 , \vrf/N198 ,
         \vrf/N197 , \vrf/N196 , \vrf/N195 , \vrf/N194 , \vrf/N193 ,
         \vrf/N192 , \vrf/N191 , \vrf/N190 , \vrf/N189 , \vrf/N188 ,
         \vrf/N187 , \vrf/N186 , \vrf/N185 , \vrf/N184 , \vrf/N183 ,
         \vrf/N182 , \vrf/N181 , \vrf/N180 , \vrf/N179 , \vrf/N178 ,
         \vrf/N177 , \vrf/N176 , \vrf/N175 , \vrf/N174 , \vrf/N173 ,
         \vrf/N172 , \vrf/N171 , \vrf/N170 , \vrf/N169 , \vrf/N168 ,
         \vrf/N167 , \vrf/N166 , \vrf/N165 , \vrf/N164 , \vrf/N163 ,
         \vrf/N162 , \vrf/N161 , \vrf/N160 , \vrf/N159 , \vrf/N158 ,
         \vrf/N157 , \vrf/N156 , \vrf/N155 , \vrf/N154 , \vrf/N153 ,
         \vrf/N152 , \vrf/N151 , \vrf/N150 , \vrf/N149 , \vrf/N148 ,
         \vrf/N147 , \vrf/N146 , \vrf/N145 , \vrf/N144 , \vrf/N143 ,
         \vrf/N142 , \vrf/N141 , \vrf/N140 , \vrf/N139 , \vrf/N138 ,
         \vrf/N137 , \vrf/N136 , \vrf/N135 , \vrf/N134 , \vrf/N133 ,
         \vrf/N132 , \vrf/N131 , \vrf/N130 , \vrf/N129 , \vrf/N128 ,
         \vrf/N127 , \vrf/N126 , \vrf/N125 , \vrf/N124 , \vrf/N123 ,
         \vrf/N122 , \vrf/N121 , \vrf/N120 , \vrf/N119 , \vrf/N118 ,
         \vrf/N116 , \vrf/N115 , \vrf/N114 , \vrf/N113 , \vrf/N112 ,
         \vrf/N111 , \vrf/N110 , \vrf/N109 , \vrf/N108 , \vrf/N107 ,
         \vrf/N106 , \vrf/N105 , \vrf/N104 , \vrf/N103 , \vrf/N102 ,
         \vrf/N101 , \vrf/N100 , \vrf/N99 , \vrf/N98 , \vrf/N97 , \vrf/N96 ,
         \vrf/N95 , \vrf/N94 , \vrf/N93 , \vrf/N92 , \vrf/N91 , \vrf/N90 ,
         \vrf/N89 , \vrf/N88 , \vrf/N87 , \vrf/N86 , \vrf/N85 , \vrf/N84 ,
         \vrf/N83 , \vrf/N82 , \vrf/N81 , \vrf/N80 , \vrf/N79 , \vrf/N78 ,
         \vrf/N77 , \vrf/N76 , \vrf/N75 , \vrf/N74 , \vrf/N73 , \vrf/N72 ,
         \vrf/N71 , \vrf/N70 , \vrf/N69 , \vrf/N68 , \vrf/N67 , \vrf/N66 ,
         \vrf/N65 , \vrf/N64 , \vrf/N63 , \vrf/N62 , \vrf/N61 , \vrf/N60 ,
         \vrf/N59 , \vrf/N58 , \vrf/N57 , \vrf/N56 , \vrf/N55 , \vrf/N54 ,
         \vrf/N53 , \vrf/N52 , \vrf/N51 , \vrf/N50 , \vrf/N49 , \vrf/N48 ,
         \vrf/N47 , \vrf/N46 , \vrf/N45 , \vrf/N44 , \vrf/N43 , \vrf/N42 ,
         \vrf/N41 , \vrf/N40 , \vrf/N39 , \vrf/N38 , \vrf/N37 , \vrf/N36 ,
         \vrf/N35 , \vrf/N34 , \vrf/N33 , \vrf/N32 , \vrf/N31 , \vrf/N30 ,
         \vrf/N29 , \vrf/N28 , \vrf/N27 , \vrf/N26 , \vrf/N25 , \vrf/N24 ,
         \vrf/N23 , \vrf/N22 , \vrf/N21 , \vrf/N20 , \vrf/N19 , \vrf/N18 ,
         \vrf/regTable[7][0] , \vrf/regTable[7][1] , \vrf/regTable[7][2] ,
         \vrf/regTable[7][3] , \vrf/regTable[7][4] , \vrf/regTable[7][5] ,
         \vrf/regTable[7][6] , \vrf/regTable[7][7] , \vrf/regTable[7][8] ,
         \vrf/regTable[7][9] , \vrf/regTable[7][10] , \vrf/regTable[7][11] ,
         \vrf/regTable[7][12] , \vrf/regTable[7][13] , \vrf/regTable[7][14] ,
         \vrf/regTable[7][15] , \vrf/regTable[7][16] , \vrf/regTable[7][17] ,
         \vrf/regTable[7][18] , \vrf/regTable[7][19] , \vrf/regTable[7][20] ,
         \vrf/regTable[7][21] , \vrf/regTable[7][22] , \vrf/regTable[7][23] ,
         \vrf/regTable[7][24] , \vrf/regTable[7][25] , \vrf/regTable[7][26] ,
         \vrf/regTable[7][27] , \vrf/regTable[7][28] , \vrf/regTable[7][29] ,
         \vrf/regTable[7][30] , \vrf/regTable[7][31] , \vrf/regTable[7][32] ,
         \vrf/regTable[7][33] , \vrf/regTable[7][34] , \vrf/regTable[7][35] ,
         \vrf/regTable[7][36] , \vrf/regTable[7][37] , \vrf/regTable[7][38] ,
         \vrf/regTable[7][39] , \vrf/regTable[7][40] , \vrf/regTable[7][41] ,
         \vrf/regTable[7][42] , \vrf/regTable[7][43] , \vrf/regTable[7][44] ,
         \vrf/regTable[7][45] , \vrf/regTable[7][46] , \vrf/regTable[7][47] ,
         \vrf/regTable[7][48] , \vrf/regTable[7][49] , \vrf/regTable[7][50] ,
         \vrf/regTable[7][51] , \vrf/regTable[7][52] , \vrf/regTable[7][53] ,
         \vrf/regTable[7][54] , \vrf/regTable[7][55] , \vrf/regTable[7][56] ,
         \vrf/regTable[7][57] , \vrf/regTable[7][58] , \vrf/regTable[7][59] ,
         \vrf/regTable[7][60] , \vrf/regTable[7][61] , \vrf/regTable[7][62] ,
         \vrf/regTable[7][63] , \vrf/regTable[7][64] , \vrf/regTable[7][65] ,
         \vrf/regTable[7][66] , \vrf/regTable[7][67] , \vrf/regTable[7][68] ,
         \vrf/regTable[7][69] , \vrf/regTable[7][70] , \vrf/regTable[7][71] ,
         \vrf/regTable[7][72] , \vrf/regTable[7][73] , \vrf/regTable[7][74] ,
         \vrf/regTable[7][75] , \vrf/regTable[7][76] , \vrf/regTable[7][77] ,
         \vrf/regTable[7][78] , \vrf/regTable[7][79] , \vrf/regTable[7][80] ,
         \vrf/regTable[7][81] , \vrf/regTable[7][82] , \vrf/regTable[7][83] ,
         \vrf/regTable[7][84] , \vrf/regTable[7][85] , \vrf/regTable[7][86] ,
         \vrf/regTable[7][87] , \vrf/regTable[7][88] , \vrf/regTable[7][89] ,
         \vrf/regTable[7][90] , \vrf/regTable[7][91] , \vrf/regTable[7][92] ,
         \vrf/regTable[7][93] , \vrf/regTable[7][94] , \vrf/regTable[7][95] ,
         \vrf/regTable[7][96] , \vrf/regTable[7][97] , \vrf/regTable[7][98] ,
         \vrf/regTable[7][99] , \vrf/regTable[7][100] , \vrf/regTable[7][101] ,
         \vrf/regTable[7][102] , \vrf/regTable[7][103] ,
         \vrf/regTable[7][104] , \vrf/regTable[7][105] ,
         \vrf/regTable[7][106] , \vrf/regTable[7][107] ,
         \vrf/regTable[7][108] , \vrf/regTable[7][109] ,
         \vrf/regTable[7][110] , \vrf/regTable[7][111] ,
         \vrf/regTable[7][112] , \vrf/regTable[7][113] ,
         \vrf/regTable[7][114] , \vrf/regTable[7][115] ,
         \vrf/regTable[7][116] , \vrf/regTable[7][117] ,
         \vrf/regTable[7][118] , \vrf/regTable[7][119] ,
         \vrf/regTable[7][120] , \vrf/regTable[7][121] ,
         \vrf/regTable[7][122] , \vrf/regTable[7][123] ,
         \vrf/regTable[7][124] , \vrf/regTable[7][125] ,
         \vrf/regTable[7][126] , \vrf/regTable[7][127] ,
         \vrf/regTable[7][128] , \vrf/regTable[7][129] ,
         \vrf/regTable[7][130] , \vrf/regTable[7][131] ,
         \vrf/regTable[7][132] , \vrf/regTable[7][133] ,
         \vrf/regTable[7][134] , \vrf/regTable[7][135] ,
         \vrf/regTable[7][136] , \vrf/regTable[7][137] ,
         \vrf/regTable[7][138] , \vrf/regTable[7][139] ,
         \vrf/regTable[7][140] , \vrf/regTable[7][141] ,
         \vrf/regTable[7][142] , \vrf/regTable[7][143] ,
         \vrf/regTable[7][144] , \vrf/regTable[7][145] ,
         \vrf/regTable[7][146] , \vrf/regTable[7][147] ,
         \vrf/regTable[7][148] , \vrf/regTable[7][149] ,
         \vrf/regTable[7][150] , \vrf/regTable[7][151] ,
         \vrf/regTable[7][152] , \vrf/regTable[7][153] ,
         \vrf/regTable[7][154] , \vrf/regTable[7][155] ,
         \vrf/regTable[7][156] , \vrf/regTable[7][157] ,
         \vrf/regTable[7][158] , \vrf/regTable[7][159] ,
         \vrf/regTable[7][160] , \vrf/regTable[7][161] ,
         \vrf/regTable[7][162] , \vrf/regTable[7][163] ,
         \vrf/regTable[7][164] , \vrf/regTable[7][165] ,
         \vrf/regTable[7][166] , \vrf/regTable[7][167] ,
         \vrf/regTable[7][168] , \vrf/regTable[7][169] ,
         \vrf/regTable[7][170] , \vrf/regTable[7][171] ,
         \vrf/regTable[7][172] , \vrf/regTable[7][173] ,
         \vrf/regTable[7][174] , \vrf/regTable[7][175] ,
         \vrf/regTable[7][176] , \vrf/regTable[7][177] ,
         \vrf/regTable[7][178] , \vrf/regTable[7][179] ,
         \vrf/regTable[7][180] , \vrf/regTable[7][181] ,
         \vrf/regTable[7][182] , \vrf/regTable[7][183] ,
         \vrf/regTable[7][184] , \vrf/regTable[7][185] ,
         \vrf/regTable[7][186] , \vrf/regTable[7][187] ,
         \vrf/regTable[7][188] , \vrf/regTable[7][189] ,
         \vrf/regTable[7][190] , \vrf/regTable[7][191] ,
         \vrf/regTable[7][192] , \vrf/regTable[7][193] ,
         \vrf/regTable[7][194] , \vrf/regTable[7][195] ,
         \vrf/regTable[7][196] , \vrf/regTable[7][197] ,
         \vrf/regTable[7][198] , \vrf/regTable[7][199] ,
         \vrf/regTable[7][200] , \vrf/regTable[7][201] ,
         \vrf/regTable[7][202] , \vrf/regTable[7][203] ,
         \vrf/regTable[7][204] , \vrf/regTable[7][205] ,
         \vrf/regTable[7][206] , \vrf/regTable[7][207] ,
         \vrf/regTable[7][208] , \vrf/regTable[7][209] ,
         \vrf/regTable[7][210] , \vrf/regTable[7][211] ,
         \vrf/regTable[7][212] , \vrf/regTable[7][213] ,
         \vrf/regTable[7][214] , \vrf/regTable[7][215] ,
         \vrf/regTable[7][216] , \vrf/regTable[7][217] ,
         \vrf/regTable[7][218] , \vrf/regTable[7][219] ,
         \vrf/regTable[7][220] , \vrf/regTable[7][221] ,
         \vrf/regTable[7][222] , \vrf/regTable[7][223] ,
         \vrf/regTable[7][224] , \vrf/regTable[7][225] ,
         \vrf/regTable[7][226] , \vrf/regTable[7][227] ,
         \vrf/regTable[7][228] , \vrf/regTable[7][229] ,
         \vrf/regTable[7][230] , \vrf/regTable[7][231] ,
         \vrf/regTable[7][232] , \vrf/regTable[7][233] ,
         \vrf/regTable[7][234] , \vrf/regTable[7][235] ,
         \vrf/regTable[7][236] , \vrf/regTable[7][237] ,
         \vrf/regTable[7][238] , \vrf/regTable[7][239] ,
         \vrf/regTable[7][240] , \vrf/regTable[7][241] ,
         \vrf/regTable[7][242] , \vrf/regTable[7][243] ,
         \vrf/regTable[7][244] , \vrf/regTable[7][245] ,
         \vrf/regTable[7][246] , \vrf/regTable[7][247] ,
         \vrf/regTable[7][248] , \vrf/regTable[7][249] ,
         \vrf/regTable[7][250] , \vrf/regTable[7][251] ,
         \vrf/regTable[7][252] , \vrf/regTable[7][253] ,
         \vrf/regTable[7][254] , \vrf/regTable[7][255] , \vrf/regTable[6][0] ,
         \vrf/regTable[6][1] , \vrf/regTable[6][2] , \vrf/regTable[6][3] ,
         \vrf/regTable[6][4] , \vrf/regTable[6][5] , \vrf/regTable[6][6] ,
         \vrf/regTable[6][7] , \vrf/regTable[6][8] , \vrf/regTable[6][9] ,
         \vrf/regTable[6][10] , \vrf/regTable[6][11] , \vrf/regTable[6][12] ,
         \vrf/regTable[6][13] , \vrf/regTable[6][14] , \vrf/regTable[6][15] ,
         \vrf/regTable[6][16] , \vrf/regTable[6][17] , \vrf/regTable[6][18] ,
         \vrf/regTable[6][19] , \vrf/regTable[6][20] , \vrf/regTable[6][21] ,
         \vrf/regTable[6][22] , \vrf/regTable[6][23] , \vrf/regTable[6][24] ,
         \vrf/regTable[6][25] , \vrf/regTable[6][26] , \vrf/regTable[6][27] ,
         \vrf/regTable[6][28] , \vrf/regTable[6][29] , \vrf/regTable[6][30] ,
         \vrf/regTable[6][31] , \vrf/regTable[6][32] , \vrf/regTable[6][33] ,
         \vrf/regTable[6][34] , \vrf/regTable[6][35] , \vrf/regTable[6][36] ,
         \vrf/regTable[6][37] , \vrf/regTable[6][38] , \vrf/regTable[6][39] ,
         \vrf/regTable[6][40] , \vrf/regTable[6][41] , \vrf/regTable[6][42] ,
         \vrf/regTable[6][43] , \vrf/regTable[6][44] , \vrf/regTable[6][45] ,
         \vrf/regTable[6][46] , \vrf/regTable[6][47] , \vrf/regTable[6][48] ,
         \vrf/regTable[6][49] , \vrf/regTable[6][50] , \vrf/regTable[6][51] ,
         \vrf/regTable[6][52] , \vrf/regTable[6][53] , \vrf/regTable[6][54] ,
         \vrf/regTable[6][55] , \vrf/regTable[6][56] , \vrf/regTable[6][57] ,
         \vrf/regTable[6][58] , \vrf/regTable[6][59] , \vrf/regTable[6][60] ,
         \vrf/regTable[6][61] , \vrf/regTable[6][62] , \vrf/regTable[6][63] ,
         \vrf/regTable[6][64] , \vrf/regTable[6][65] , \vrf/regTable[6][66] ,
         \vrf/regTable[6][67] , \vrf/regTable[6][68] , \vrf/regTable[6][69] ,
         \vrf/regTable[6][70] , \vrf/regTable[6][71] , \vrf/regTable[6][72] ,
         \vrf/regTable[6][73] , \vrf/regTable[6][74] , \vrf/regTable[6][75] ,
         \vrf/regTable[6][76] , \vrf/regTable[6][77] , \vrf/regTable[6][78] ,
         \vrf/regTable[6][79] , \vrf/regTable[6][80] , \vrf/regTable[6][81] ,
         \vrf/regTable[6][82] , \vrf/regTable[6][83] , \vrf/regTable[6][84] ,
         \vrf/regTable[6][85] , \vrf/regTable[6][86] , \vrf/regTable[6][87] ,
         \vrf/regTable[6][88] , \vrf/regTable[6][89] , \vrf/regTable[6][90] ,
         \vrf/regTable[6][91] , \vrf/regTable[6][92] , \vrf/regTable[6][93] ,
         \vrf/regTable[6][94] , \vrf/regTable[6][95] , \vrf/regTable[6][96] ,
         \vrf/regTable[6][97] , \vrf/regTable[6][98] , \vrf/regTable[6][99] ,
         \vrf/regTable[6][100] , \vrf/regTable[6][101] ,
         \vrf/regTable[6][102] , \vrf/regTable[6][103] ,
         \vrf/regTable[6][104] , \vrf/regTable[6][105] ,
         \vrf/regTable[6][106] , \vrf/regTable[6][107] ,
         \vrf/regTable[6][108] , \vrf/regTable[6][109] ,
         \vrf/regTable[6][110] , \vrf/regTable[6][111] ,
         \vrf/regTable[6][112] , \vrf/regTable[6][113] ,
         \vrf/regTable[6][114] , \vrf/regTable[6][115] ,
         \vrf/regTable[6][116] , \vrf/regTable[6][117] ,
         \vrf/regTable[6][118] , \vrf/regTable[6][119] ,
         \vrf/regTable[6][120] , \vrf/regTable[6][121] ,
         \vrf/regTable[6][122] , \vrf/regTable[6][123] ,
         \vrf/regTable[6][124] , \vrf/regTable[6][125] ,
         \vrf/regTable[6][126] , \vrf/regTable[6][127] ,
         \vrf/regTable[6][128] , \vrf/regTable[6][129] ,
         \vrf/regTable[6][130] , \vrf/regTable[6][131] ,
         \vrf/regTable[6][132] , \vrf/regTable[6][133] ,
         \vrf/regTable[6][134] , \vrf/regTable[6][135] ,
         \vrf/regTable[6][136] , \vrf/regTable[6][137] ,
         \vrf/regTable[6][138] , \vrf/regTable[6][139] ,
         \vrf/regTable[6][140] , \vrf/regTable[6][141] ,
         \vrf/regTable[6][142] , \vrf/regTable[6][143] ,
         \vrf/regTable[6][144] , \vrf/regTable[6][145] ,
         \vrf/regTable[6][146] , \vrf/regTable[6][147] ,
         \vrf/regTable[6][148] , \vrf/regTable[6][149] ,
         \vrf/regTable[6][150] , \vrf/regTable[6][151] ,
         \vrf/regTable[6][152] , \vrf/regTable[6][153] ,
         \vrf/regTable[6][154] , \vrf/regTable[6][155] ,
         \vrf/regTable[6][156] , \vrf/regTable[6][157] ,
         \vrf/regTable[6][158] , \vrf/regTable[6][159] ,
         \vrf/regTable[6][160] , \vrf/regTable[6][161] ,
         \vrf/regTable[6][162] , \vrf/regTable[6][163] ,
         \vrf/regTable[6][164] , \vrf/regTable[6][165] ,
         \vrf/regTable[6][166] , \vrf/regTable[6][167] ,
         \vrf/regTable[6][168] , \vrf/regTable[6][169] ,
         \vrf/regTable[6][170] , \vrf/regTable[6][171] ,
         \vrf/regTable[6][172] , \vrf/regTable[6][173] ,
         \vrf/regTable[6][174] , \vrf/regTable[6][175] ,
         \vrf/regTable[6][176] , \vrf/regTable[6][177] ,
         \vrf/regTable[6][178] , \vrf/regTable[6][179] ,
         \vrf/regTable[6][180] , \vrf/regTable[6][181] ,
         \vrf/regTable[6][182] , \vrf/regTable[6][183] ,
         \vrf/regTable[6][184] , \vrf/regTable[6][185] ,
         \vrf/regTable[6][186] , \vrf/regTable[6][187] ,
         \vrf/regTable[6][188] , \vrf/regTable[6][189] ,
         \vrf/regTable[6][190] , \vrf/regTable[6][191] ,
         \vrf/regTable[6][192] , \vrf/regTable[6][193] ,
         \vrf/regTable[6][194] , \vrf/regTable[6][195] ,
         \vrf/regTable[6][196] , \vrf/regTable[6][197] ,
         \vrf/regTable[6][198] , \vrf/regTable[6][199] ,
         \vrf/regTable[6][200] , \vrf/regTable[6][201] ,
         \vrf/regTable[6][202] , \vrf/regTable[6][203] ,
         \vrf/regTable[6][204] , \vrf/regTable[6][205] ,
         \vrf/regTable[6][206] , \vrf/regTable[6][207] ,
         \vrf/regTable[6][208] , \vrf/regTable[6][209] ,
         \vrf/regTable[6][210] , \vrf/regTable[6][211] ,
         \vrf/regTable[6][212] , \vrf/regTable[6][213] ,
         \vrf/regTable[6][214] , \vrf/regTable[6][215] ,
         \vrf/regTable[6][216] , \vrf/regTable[6][217] ,
         \vrf/regTable[6][218] , \vrf/regTable[6][219] ,
         \vrf/regTable[6][220] , \vrf/regTable[6][221] ,
         \vrf/regTable[6][222] , \vrf/regTable[6][223] ,
         \vrf/regTable[6][224] , \vrf/regTable[6][225] ,
         \vrf/regTable[6][226] , \vrf/regTable[6][227] ,
         \vrf/regTable[6][228] , \vrf/regTable[6][229] ,
         \vrf/regTable[6][230] , \vrf/regTable[6][231] ,
         \vrf/regTable[6][232] , \vrf/regTable[6][233] ,
         \vrf/regTable[6][234] , \vrf/regTable[6][235] ,
         \vrf/regTable[6][236] , \vrf/regTable[6][237] ,
         \vrf/regTable[6][238] , \vrf/regTable[6][239] ,
         \vrf/regTable[6][240] , \vrf/regTable[6][241] ,
         \vrf/regTable[6][242] , \vrf/regTable[6][243] ,
         \vrf/regTable[6][244] , \vrf/regTable[6][245] ,
         \vrf/regTable[6][246] , \vrf/regTable[6][247] ,
         \vrf/regTable[6][248] , \vrf/regTable[6][249] ,
         \vrf/regTable[6][250] , \vrf/regTable[6][251] ,
         \vrf/regTable[6][252] , \vrf/regTable[6][253] ,
         \vrf/regTable[6][254] , \vrf/regTable[6][255] , \vrf/regTable[5][0] ,
         \vrf/regTable[5][1] , \vrf/regTable[5][2] , \vrf/regTable[5][3] ,
         \vrf/regTable[5][4] , \vrf/regTable[5][5] , \vrf/regTable[5][6] ,
         \vrf/regTable[5][7] , \vrf/regTable[5][8] , \vrf/regTable[5][9] ,
         \vrf/regTable[5][10] , \vrf/regTable[5][11] , \vrf/regTable[5][12] ,
         \vrf/regTable[5][13] , \vrf/regTable[5][14] , \vrf/regTable[5][15] ,
         \vrf/regTable[5][16] , \vrf/regTable[5][17] , \vrf/regTable[5][18] ,
         \vrf/regTable[5][19] , \vrf/regTable[5][20] , \vrf/regTable[5][21] ,
         \vrf/regTable[5][22] , \vrf/regTable[5][23] , \vrf/regTable[5][24] ,
         \vrf/regTable[5][25] , \vrf/regTable[5][26] , \vrf/regTable[5][27] ,
         \vrf/regTable[5][28] , \vrf/regTable[5][29] , \vrf/regTable[5][30] ,
         \vrf/regTable[5][31] , \vrf/regTable[5][32] , \vrf/regTable[5][33] ,
         \vrf/regTable[5][34] , \vrf/regTable[5][35] , \vrf/regTable[5][36] ,
         \vrf/regTable[5][37] , \vrf/regTable[5][38] , \vrf/regTable[5][39] ,
         \vrf/regTable[5][40] , \vrf/regTable[5][41] , \vrf/regTable[5][42] ,
         \vrf/regTable[5][43] , \vrf/regTable[5][44] , \vrf/regTable[5][45] ,
         \vrf/regTable[5][46] , \vrf/regTable[5][47] , \vrf/regTable[5][48] ,
         \vrf/regTable[5][49] , \vrf/regTable[5][50] , \vrf/regTable[5][51] ,
         \vrf/regTable[5][52] , \vrf/regTable[5][53] , \vrf/regTable[5][54] ,
         \vrf/regTable[5][55] , \vrf/regTable[5][56] , \vrf/regTable[5][57] ,
         \vrf/regTable[5][58] , \vrf/regTable[5][59] , \vrf/regTable[5][60] ,
         \vrf/regTable[5][61] , \vrf/regTable[5][62] , \vrf/regTable[5][63] ,
         \vrf/regTable[5][64] , \vrf/regTable[5][65] , \vrf/regTable[5][66] ,
         \vrf/regTable[5][67] , \vrf/regTable[5][68] , \vrf/regTable[5][69] ,
         \vrf/regTable[5][70] , \vrf/regTable[5][71] , \vrf/regTable[5][72] ,
         \vrf/regTable[5][73] , \vrf/regTable[5][74] , \vrf/regTable[5][75] ,
         \vrf/regTable[5][76] , \vrf/regTable[5][77] , \vrf/regTable[5][78] ,
         \vrf/regTable[5][79] , \vrf/regTable[5][80] , \vrf/regTable[5][81] ,
         \vrf/regTable[5][82] , \vrf/regTable[5][83] , \vrf/regTable[5][84] ,
         \vrf/regTable[5][85] , \vrf/regTable[5][86] , \vrf/regTable[5][87] ,
         \vrf/regTable[5][88] , \vrf/regTable[5][89] , \vrf/regTable[5][90] ,
         \vrf/regTable[5][91] , \vrf/regTable[5][92] , \vrf/regTable[5][93] ,
         \vrf/regTable[5][94] , \vrf/regTable[5][95] , \vrf/regTable[5][96] ,
         \vrf/regTable[5][97] , \vrf/regTable[5][98] , \vrf/regTable[5][99] ,
         \vrf/regTable[5][100] , \vrf/regTable[5][101] ,
         \vrf/regTable[5][102] , \vrf/regTable[5][103] ,
         \vrf/regTable[5][104] , \vrf/regTable[5][105] ,
         \vrf/regTable[5][106] , \vrf/regTable[5][107] ,
         \vrf/regTable[5][108] , \vrf/regTable[5][109] ,
         \vrf/regTable[5][110] , \vrf/regTable[5][111] ,
         \vrf/regTable[5][112] , \vrf/regTable[5][113] ,
         \vrf/regTable[5][114] , \vrf/regTable[5][115] ,
         \vrf/regTable[5][116] , \vrf/regTable[5][117] ,
         \vrf/regTable[5][118] , \vrf/regTable[5][119] ,
         \vrf/regTable[5][120] , \vrf/regTable[5][121] ,
         \vrf/regTable[5][122] , \vrf/regTable[5][123] ,
         \vrf/regTable[5][124] , \vrf/regTable[5][125] ,
         \vrf/regTable[5][126] , \vrf/regTable[5][127] ,
         \vrf/regTable[5][128] , \vrf/regTable[5][129] ,
         \vrf/regTable[5][130] , \vrf/regTable[5][131] ,
         \vrf/regTable[5][132] , \vrf/regTable[5][133] ,
         \vrf/regTable[5][134] , \vrf/regTable[5][135] ,
         \vrf/regTable[5][136] , \vrf/regTable[5][137] ,
         \vrf/regTable[5][138] , \vrf/regTable[5][139] ,
         \vrf/regTable[5][140] , \vrf/regTable[5][141] ,
         \vrf/regTable[5][142] , \vrf/regTable[5][143] ,
         \vrf/regTable[5][144] , \vrf/regTable[5][145] ,
         \vrf/regTable[5][146] , \vrf/regTable[5][147] ,
         \vrf/regTable[5][148] , \vrf/regTable[5][149] ,
         \vrf/regTable[5][150] , \vrf/regTable[5][151] ,
         \vrf/regTable[5][152] , \vrf/regTable[5][153] ,
         \vrf/regTable[5][154] , \vrf/regTable[5][155] ,
         \vrf/regTable[5][156] , \vrf/regTable[5][157] ,
         \vrf/regTable[5][158] , \vrf/regTable[5][159] ,
         \vrf/regTable[5][160] , \vrf/regTable[5][161] ,
         \vrf/regTable[5][162] , \vrf/regTable[5][163] ,
         \vrf/regTable[5][164] , \vrf/regTable[5][165] ,
         \vrf/regTable[5][166] , \vrf/regTable[5][167] ,
         \vrf/regTable[5][168] , \vrf/regTable[5][169] ,
         \vrf/regTable[5][170] , \vrf/regTable[5][171] ,
         \vrf/regTable[5][172] , \vrf/regTable[5][173] ,
         \vrf/regTable[5][174] , \vrf/regTable[5][175] ,
         \vrf/regTable[5][176] , \vrf/regTable[5][177] ,
         \vrf/regTable[5][178] , \vrf/regTable[5][179] ,
         \vrf/regTable[5][180] , \vrf/regTable[5][181] ,
         \vrf/regTable[5][182] , \vrf/regTable[5][183] ,
         \vrf/regTable[5][184] , \vrf/regTable[5][185] ,
         \vrf/regTable[5][186] , \vrf/regTable[5][187] ,
         \vrf/regTable[5][188] , \vrf/regTable[5][189] ,
         \vrf/regTable[5][190] , \vrf/regTable[5][191] ,
         \vrf/regTable[5][192] , \vrf/regTable[5][193] ,
         \vrf/regTable[5][194] , \vrf/regTable[5][195] ,
         \vrf/regTable[5][196] , \vrf/regTable[5][197] ,
         \vrf/regTable[5][198] , \vrf/regTable[5][199] ,
         \vrf/regTable[5][200] , \vrf/regTable[5][201] ,
         \vrf/regTable[5][202] , \vrf/regTable[5][203] ,
         \vrf/regTable[5][204] , \vrf/regTable[5][205] ,
         \vrf/regTable[5][206] , \vrf/regTable[5][207] ,
         \vrf/regTable[5][208] , \vrf/regTable[5][209] ,
         \vrf/regTable[5][210] , \vrf/regTable[5][211] ,
         \vrf/regTable[5][212] , \vrf/regTable[5][213] ,
         \vrf/regTable[5][214] , \vrf/regTable[5][215] ,
         \vrf/regTable[5][216] , \vrf/regTable[5][217] ,
         \vrf/regTable[5][218] , \vrf/regTable[5][219] ,
         \vrf/regTable[5][220] , \vrf/regTable[5][221] ,
         \vrf/regTable[5][222] , \vrf/regTable[5][223] ,
         \vrf/regTable[5][224] , \vrf/regTable[5][225] ,
         \vrf/regTable[5][226] , \vrf/regTable[5][227] ,
         \vrf/regTable[5][228] , \vrf/regTable[5][229] ,
         \vrf/regTable[5][230] , \vrf/regTable[5][231] ,
         \vrf/regTable[5][232] , \vrf/regTable[5][233] ,
         \vrf/regTable[5][234] , \vrf/regTable[5][235] ,
         \vrf/regTable[5][236] , \vrf/regTable[5][237] ,
         \vrf/regTable[5][238] , \vrf/regTable[5][239] ,
         \vrf/regTable[5][240] , \vrf/regTable[5][241] ,
         \vrf/regTable[5][242] , \vrf/regTable[5][243] ,
         \vrf/regTable[5][244] , \vrf/regTable[5][245] ,
         \vrf/regTable[5][246] , \vrf/regTable[5][247] ,
         \vrf/regTable[5][248] , \vrf/regTable[5][249] ,
         \vrf/regTable[5][250] , \vrf/regTable[5][251] ,
         \vrf/regTable[5][252] , \vrf/regTable[5][253] ,
         \vrf/regTable[5][254] , \vrf/regTable[5][255] , \vrf/regTable[4][0] ,
         \vrf/regTable[4][1] , \vrf/regTable[4][2] , \vrf/regTable[4][3] ,
         \vrf/regTable[4][4] , \vrf/regTable[4][5] , \vrf/regTable[4][6] ,
         \vrf/regTable[4][7] , \vrf/regTable[4][8] , \vrf/regTable[4][9] ,
         \vrf/regTable[4][10] , \vrf/regTable[4][11] , \vrf/regTable[4][12] ,
         \vrf/regTable[4][13] , \vrf/regTable[4][14] , \vrf/regTable[4][15] ,
         \vrf/regTable[4][16] , \vrf/regTable[4][17] , \vrf/regTable[4][18] ,
         \vrf/regTable[4][19] , \vrf/regTable[4][20] , \vrf/regTable[4][21] ,
         \vrf/regTable[4][22] , \vrf/regTable[4][23] , \vrf/regTable[4][24] ,
         \vrf/regTable[4][25] , \vrf/regTable[4][26] , \vrf/regTable[4][27] ,
         \vrf/regTable[4][28] , \vrf/regTable[4][29] , \vrf/regTable[4][30] ,
         \vrf/regTable[4][31] , \vrf/regTable[4][32] , \vrf/regTable[4][33] ,
         \vrf/regTable[4][34] , \vrf/regTable[4][35] , \vrf/regTable[4][36] ,
         \vrf/regTable[4][37] , \vrf/regTable[4][38] , \vrf/regTable[4][39] ,
         \vrf/regTable[4][40] , \vrf/regTable[4][41] , \vrf/regTable[4][42] ,
         \vrf/regTable[4][43] , \vrf/regTable[4][44] , \vrf/regTable[4][45] ,
         \vrf/regTable[4][46] , \vrf/regTable[4][47] , \vrf/regTable[4][48] ,
         \vrf/regTable[4][49] , \vrf/regTable[4][50] , \vrf/regTable[4][51] ,
         \vrf/regTable[4][52] , \vrf/regTable[4][53] , \vrf/regTable[4][54] ,
         \vrf/regTable[4][55] , \vrf/regTable[4][56] , \vrf/regTable[4][57] ,
         \vrf/regTable[4][58] , \vrf/regTable[4][59] , \vrf/regTable[4][60] ,
         \vrf/regTable[4][61] , \vrf/regTable[4][62] , \vrf/regTable[4][63] ,
         \vrf/regTable[4][64] , \vrf/regTable[4][65] , \vrf/regTable[4][66] ,
         \vrf/regTable[4][67] , \vrf/regTable[4][68] , \vrf/regTable[4][69] ,
         \vrf/regTable[4][70] , \vrf/regTable[4][71] , \vrf/regTable[4][72] ,
         \vrf/regTable[4][73] , \vrf/regTable[4][74] , \vrf/regTable[4][75] ,
         \vrf/regTable[4][76] , \vrf/regTable[4][77] , \vrf/regTable[4][78] ,
         \vrf/regTable[4][79] , \vrf/regTable[4][80] , \vrf/regTable[4][81] ,
         \vrf/regTable[4][82] , \vrf/regTable[4][83] , \vrf/regTable[4][84] ,
         \vrf/regTable[4][85] , \vrf/regTable[4][86] , \vrf/regTable[4][87] ,
         \vrf/regTable[4][88] , \vrf/regTable[4][89] , \vrf/regTable[4][90] ,
         \vrf/regTable[4][91] , \vrf/regTable[4][92] , \vrf/regTable[4][93] ,
         \vrf/regTable[4][94] , \vrf/regTable[4][95] , \vrf/regTable[4][96] ,
         \vrf/regTable[4][97] , \vrf/regTable[4][98] , \vrf/regTable[4][99] ,
         \vrf/regTable[4][100] , \vrf/regTable[4][101] ,
         \vrf/regTable[4][102] , \vrf/regTable[4][103] ,
         \vrf/regTable[4][104] , \vrf/regTable[4][105] ,
         \vrf/regTable[4][106] , \vrf/regTable[4][107] ,
         \vrf/regTable[4][108] , \vrf/regTable[4][109] ,
         \vrf/regTable[4][110] , \vrf/regTable[4][111] ,
         \vrf/regTable[4][112] , \vrf/regTable[4][113] ,
         \vrf/regTable[4][114] , \vrf/regTable[4][115] ,
         \vrf/regTable[4][116] , \vrf/regTable[4][117] ,
         \vrf/regTable[4][118] , \vrf/regTable[4][119] ,
         \vrf/regTable[4][120] , \vrf/regTable[4][121] ,
         \vrf/regTable[4][122] , \vrf/regTable[4][123] ,
         \vrf/regTable[4][124] , \vrf/regTable[4][125] ,
         \vrf/regTable[4][126] , \vrf/regTable[4][127] ,
         \vrf/regTable[4][128] , \vrf/regTable[4][129] ,
         \vrf/regTable[4][130] , \vrf/regTable[4][131] ,
         \vrf/regTable[4][132] , \vrf/regTable[4][133] ,
         \vrf/regTable[4][134] , \vrf/regTable[4][135] ,
         \vrf/regTable[4][136] , \vrf/regTable[4][137] ,
         \vrf/regTable[4][138] , \vrf/regTable[4][139] ,
         \vrf/regTable[4][140] , \vrf/regTable[4][141] ,
         \vrf/regTable[4][142] , \vrf/regTable[4][143] ,
         \vrf/regTable[4][144] , \vrf/regTable[4][145] ,
         \vrf/regTable[4][146] , \vrf/regTable[4][147] ,
         \vrf/regTable[4][148] , \vrf/regTable[4][149] ,
         \vrf/regTable[4][150] , \vrf/regTable[4][151] ,
         \vrf/regTable[4][152] , \vrf/regTable[4][153] ,
         \vrf/regTable[4][154] , \vrf/regTable[4][155] ,
         \vrf/regTable[4][156] , \vrf/regTable[4][157] ,
         \vrf/regTable[4][158] , \vrf/regTable[4][159] ,
         \vrf/regTable[4][160] , \vrf/regTable[4][161] ,
         \vrf/regTable[4][162] , \vrf/regTable[4][163] ,
         \vrf/regTable[4][164] , \vrf/regTable[4][165] ,
         \vrf/regTable[4][166] , \vrf/regTable[4][167] ,
         \vrf/regTable[4][168] , \vrf/regTable[4][169] ,
         \vrf/regTable[4][170] , \vrf/regTable[4][171] ,
         \vrf/regTable[4][172] , \vrf/regTable[4][173] ,
         \vrf/regTable[4][174] , \vrf/regTable[4][175] ,
         \vrf/regTable[4][176] , \vrf/regTable[4][177] ,
         \vrf/regTable[4][178] , \vrf/regTable[4][179] ,
         \vrf/regTable[4][180] , \vrf/regTable[4][181] ,
         \vrf/regTable[4][182] , \vrf/regTable[4][183] ,
         \vrf/regTable[4][184] , \vrf/regTable[4][185] ,
         \vrf/regTable[4][186] , \vrf/regTable[4][187] ,
         \vrf/regTable[4][188] , \vrf/regTable[4][189] ,
         \vrf/regTable[4][190] , \vrf/regTable[4][191] ,
         \vrf/regTable[4][192] , \vrf/regTable[4][193] ,
         \vrf/regTable[4][194] , \vrf/regTable[4][195] ,
         \vrf/regTable[4][196] , \vrf/regTable[4][197] ,
         \vrf/regTable[4][198] , \vrf/regTable[4][199] ,
         \vrf/regTable[4][200] , \vrf/regTable[4][201] ,
         \vrf/regTable[4][202] , \vrf/regTable[4][203] ,
         \vrf/regTable[4][204] , \vrf/regTable[4][205] ,
         \vrf/regTable[4][206] , \vrf/regTable[4][207] ,
         \vrf/regTable[4][208] , \vrf/regTable[4][209] ,
         \vrf/regTable[4][210] , \vrf/regTable[4][211] ,
         \vrf/regTable[4][212] , \vrf/regTable[4][213] ,
         \vrf/regTable[4][214] , \vrf/regTable[4][215] ,
         \vrf/regTable[4][216] , \vrf/regTable[4][217] ,
         \vrf/regTable[4][218] , \vrf/regTable[4][219] ,
         \vrf/regTable[4][220] , \vrf/regTable[4][221] ,
         \vrf/regTable[4][222] , \vrf/regTable[4][223] ,
         \vrf/regTable[4][224] , \vrf/regTable[4][225] ,
         \vrf/regTable[4][226] , \vrf/regTable[4][227] ,
         \vrf/regTable[4][228] , \vrf/regTable[4][229] ,
         \vrf/regTable[4][230] , \vrf/regTable[4][231] ,
         \vrf/regTable[4][232] , \vrf/regTable[4][233] ,
         \vrf/regTable[4][234] , \vrf/regTable[4][235] ,
         \vrf/regTable[4][236] , \vrf/regTable[4][237] ,
         \vrf/regTable[4][238] , \vrf/regTable[4][239] ,
         \vrf/regTable[4][240] , \vrf/regTable[4][241] ,
         \vrf/regTable[4][242] , \vrf/regTable[4][243] ,
         \vrf/regTable[4][244] , \vrf/regTable[4][245] ,
         \vrf/regTable[4][246] , \vrf/regTable[4][247] ,
         \vrf/regTable[4][248] , \vrf/regTable[4][249] ,
         \vrf/regTable[4][250] , \vrf/regTable[4][251] ,
         \vrf/regTable[4][252] , \vrf/regTable[4][253] ,
         \vrf/regTable[4][254] , \vrf/regTable[4][255] , \vrf/regTable[3][0] ,
         \vrf/regTable[3][1] , \vrf/regTable[3][2] , \vrf/regTable[3][3] ,
         \vrf/regTable[3][4] , \vrf/regTable[3][5] , \vrf/regTable[3][6] ,
         \vrf/regTable[3][7] , \vrf/regTable[3][8] , \vrf/regTable[3][9] ,
         \vrf/regTable[3][10] , \vrf/regTable[3][11] , \vrf/regTable[3][12] ,
         \vrf/regTable[3][13] , \vrf/regTable[3][14] , \vrf/regTable[3][15] ,
         \vrf/regTable[3][16] , \vrf/regTable[3][17] , \vrf/regTable[3][18] ,
         \vrf/regTable[3][19] , \vrf/regTable[3][20] , \vrf/regTable[3][21] ,
         \vrf/regTable[3][22] , \vrf/regTable[3][23] , \vrf/regTable[3][24] ,
         \vrf/regTable[3][25] , \vrf/regTable[3][26] , \vrf/regTable[3][27] ,
         \vrf/regTable[3][28] , \vrf/regTable[3][29] , \vrf/regTable[3][30] ,
         \vrf/regTable[3][31] , \vrf/regTable[3][32] , \vrf/regTable[3][33] ,
         \vrf/regTable[3][34] , \vrf/regTable[3][35] , \vrf/regTable[3][36] ,
         \vrf/regTable[3][37] , \vrf/regTable[3][38] , \vrf/regTable[3][39] ,
         \vrf/regTable[3][40] , \vrf/regTable[3][41] , \vrf/regTable[3][42] ,
         \vrf/regTable[3][43] , \vrf/regTable[3][44] , \vrf/regTable[3][45] ,
         \vrf/regTable[3][46] , \vrf/regTable[3][47] , \vrf/regTable[3][48] ,
         \vrf/regTable[3][49] , \vrf/regTable[3][50] , \vrf/regTable[3][51] ,
         \vrf/regTable[3][52] , \vrf/regTable[3][53] , \vrf/regTable[3][54] ,
         \vrf/regTable[3][55] , \vrf/regTable[3][56] , \vrf/regTable[3][57] ,
         \vrf/regTable[3][58] , \vrf/regTable[3][59] , \vrf/regTable[3][60] ,
         \vrf/regTable[3][61] , \vrf/regTable[3][62] , \vrf/regTable[3][63] ,
         \vrf/regTable[3][64] , \vrf/regTable[3][65] , \vrf/regTable[3][66] ,
         \vrf/regTable[3][67] , \vrf/regTable[3][68] , \vrf/regTable[3][69] ,
         \vrf/regTable[3][70] , \vrf/regTable[3][71] , \vrf/regTable[3][72] ,
         \vrf/regTable[3][73] , \vrf/regTable[3][74] , \vrf/regTable[3][75] ,
         \vrf/regTable[3][76] , \vrf/regTable[3][77] , \vrf/regTable[3][78] ,
         \vrf/regTable[3][79] , \vrf/regTable[3][80] , \vrf/regTable[3][81] ,
         \vrf/regTable[3][82] , \vrf/regTable[3][83] , \vrf/regTable[3][84] ,
         \vrf/regTable[3][85] , \vrf/regTable[3][86] , \vrf/regTable[3][87] ,
         \vrf/regTable[3][88] , \vrf/regTable[3][89] , \vrf/regTable[3][90] ,
         \vrf/regTable[3][91] , \vrf/regTable[3][92] , \vrf/regTable[3][93] ,
         \vrf/regTable[3][94] , \vrf/regTable[3][95] , \vrf/regTable[3][96] ,
         \vrf/regTable[3][97] , \vrf/regTable[3][98] , \vrf/regTable[3][99] ,
         \vrf/regTable[3][100] , \vrf/regTable[3][101] ,
         \vrf/regTable[3][102] , \vrf/regTable[3][103] ,
         \vrf/regTable[3][104] , \vrf/regTable[3][105] ,
         \vrf/regTable[3][106] , \vrf/regTable[3][107] ,
         \vrf/regTable[3][108] , \vrf/regTable[3][109] ,
         \vrf/regTable[3][110] , \vrf/regTable[3][111] ,
         \vrf/regTable[3][112] , \vrf/regTable[3][113] ,
         \vrf/regTable[3][114] , \vrf/regTable[3][115] ,
         \vrf/regTable[3][116] , \vrf/regTable[3][117] ,
         \vrf/regTable[3][118] , \vrf/regTable[3][119] ,
         \vrf/regTable[3][120] , \vrf/regTable[3][121] ,
         \vrf/regTable[3][122] , \vrf/regTable[3][123] ,
         \vrf/regTable[3][124] , \vrf/regTable[3][125] ,
         \vrf/regTable[3][126] , \vrf/regTable[3][127] ,
         \vrf/regTable[3][128] , \vrf/regTable[3][129] ,
         \vrf/regTable[3][130] , \vrf/regTable[3][131] ,
         \vrf/regTable[3][132] , \vrf/regTable[3][133] ,
         \vrf/regTable[3][134] , \vrf/regTable[3][135] ,
         \vrf/regTable[3][136] , \vrf/regTable[3][137] ,
         \vrf/regTable[3][138] , \vrf/regTable[3][139] ,
         \vrf/regTable[3][140] , \vrf/regTable[3][141] ,
         \vrf/regTable[3][142] , \vrf/regTable[3][143] ,
         \vrf/regTable[3][144] , \vrf/regTable[3][145] ,
         \vrf/regTable[3][146] , \vrf/regTable[3][147] ,
         \vrf/regTable[3][148] , \vrf/regTable[3][149] ,
         \vrf/regTable[3][150] , \vrf/regTable[3][151] ,
         \vrf/regTable[3][152] , \vrf/regTable[3][153] ,
         \vrf/regTable[3][154] , \vrf/regTable[3][155] ,
         \vrf/regTable[3][156] , \vrf/regTable[3][157] ,
         \vrf/regTable[3][158] , \vrf/regTable[3][159] ,
         \vrf/regTable[3][160] , \vrf/regTable[3][161] ,
         \vrf/regTable[3][162] , \vrf/regTable[3][163] ,
         \vrf/regTable[3][164] , \vrf/regTable[3][165] ,
         \vrf/regTable[3][166] , \vrf/regTable[3][167] ,
         \vrf/regTable[3][168] , \vrf/regTable[3][169] ,
         \vrf/regTable[3][170] , \vrf/regTable[3][171] ,
         \vrf/regTable[3][172] , \vrf/regTable[3][173] ,
         \vrf/regTable[3][174] , \vrf/regTable[3][175] ,
         \vrf/regTable[3][176] , \vrf/regTable[3][177] ,
         \vrf/regTable[3][178] , \vrf/regTable[3][179] ,
         \vrf/regTable[3][180] , \vrf/regTable[3][181] ,
         \vrf/regTable[3][182] , \vrf/regTable[3][183] ,
         \vrf/regTable[3][184] , \vrf/regTable[3][185] ,
         \vrf/regTable[3][186] , \vrf/regTable[3][187] ,
         \vrf/regTable[3][188] , \vrf/regTable[3][189] ,
         \vrf/regTable[3][190] , \vrf/regTable[3][191] ,
         \vrf/regTable[3][192] , \vrf/regTable[3][193] ,
         \vrf/regTable[3][194] , \vrf/regTable[3][195] ,
         \vrf/regTable[3][196] , \vrf/regTable[3][197] ,
         \vrf/regTable[3][198] , \vrf/regTable[3][199] ,
         \vrf/regTable[3][200] , \vrf/regTable[3][201] ,
         \vrf/regTable[3][202] , \vrf/regTable[3][203] ,
         \vrf/regTable[3][204] , \vrf/regTable[3][205] ,
         \vrf/regTable[3][206] , \vrf/regTable[3][207] ,
         \vrf/regTable[3][208] , \vrf/regTable[3][209] ,
         \vrf/regTable[3][210] , \vrf/regTable[3][211] ,
         \vrf/regTable[3][212] , \vrf/regTable[3][213] ,
         \vrf/regTable[3][214] , \vrf/regTable[3][215] ,
         \vrf/regTable[3][216] , \vrf/regTable[3][217] ,
         \vrf/regTable[3][218] , \vrf/regTable[3][219] ,
         \vrf/regTable[3][220] , \vrf/regTable[3][221] ,
         \vrf/regTable[3][222] , \vrf/regTable[3][223] ,
         \vrf/regTable[3][224] , \vrf/regTable[3][225] ,
         \vrf/regTable[3][226] , \vrf/regTable[3][227] ,
         \vrf/regTable[3][228] , \vrf/regTable[3][229] ,
         \vrf/regTable[3][230] , \vrf/regTable[3][231] ,
         \vrf/regTable[3][232] , \vrf/regTable[3][233] ,
         \vrf/regTable[3][234] , \vrf/regTable[3][235] ,
         \vrf/regTable[3][236] , \vrf/regTable[3][237] ,
         \vrf/regTable[3][238] , \vrf/regTable[3][239] ,
         \vrf/regTable[3][240] , \vrf/regTable[3][241] ,
         \vrf/regTable[3][242] , \vrf/regTable[3][243] ,
         \vrf/regTable[3][244] , \vrf/regTable[3][245] ,
         \vrf/regTable[3][246] , \vrf/regTable[3][247] ,
         \vrf/regTable[3][248] , \vrf/regTable[3][249] ,
         \vrf/regTable[3][250] , \vrf/regTable[3][251] ,
         \vrf/regTable[3][252] , \vrf/regTable[3][253] ,
         \vrf/regTable[3][254] , \vrf/regTable[3][255] , \vrf/regTable[2][0] ,
         \vrf/regTable[2][1] , \vrf/regTable[2][2] , \vrf/regTable[2][3] ,
         \vrf/regTable[2][4] , \vrf/regTable[2][5] , \vrf/regTable[2][6] ,
         \vrf/regTable[2][7] , \vrf/regTable[2][8] , \vrf/regTable[2][9] ,
         \vrf/regTable[2][10] , \vrf/regTable[2][11] , \vrf/regTable[2][12] ,
         \vrf/regTable[2][13] , \vrf/regTable[2][14] , \vrf/regTable[2][15] ,
         \vrf/regTable[2][16] , \vrf/regTable[2][17] , \vrf/regTable[2][18] ,
         \vrf/regTable[2][19] , \vrf/regTable[2][20] , \vrf/regTable[2][21] ,
         \vrf/regTable[2][22] , \vrf/regTable[2][23] , \vrf/regTable[2][24] ,
         \vrf/regTable[2][25] , \vrf/regTable[2][26] , \vrf/regTable[2][27] ,
         \vrf/regTable[2][28] , \vrf/regTable[2][29] , \vrf/regTable[2][30] ,
         \vrf/regTable[2][31] , \vrf/regTable[2][32] , \vrf/regTable[2][33] ,
         \vrf/regTable[2][34] , \vrf/regTable[2][35] , \vrf/regTable[2][36] ,
         \vrf/regTable[2][37] , \vrf/regTable[2][38] , \vrf/regTable[2][39] ,
         \vrf/regTable[2][40] , \vrf/regTable[2][41] , \vrf/regTable[2][42] ,
         \vrf/regTable[2][43] , \vrf/regTable[2][44] , \vrf/regTable[2][45] ,
         \vrf/regTable[2][46] , \vrf/regTable[2][47] , \vrf/regTable[2][48] ,
         \vrf/regTable[2][49] , \vrf/regTable[2][50] , \vrf/regTable[2][51] ,
         \vrf/regTable[2][52] , \vrf/regTable[2][53] , \vrf/regTable[2][54] ,
         \vrf/regTable[2][55] , \vrf/regTable[2][56] , \vrf/regTable[2][57] ,
         \vrf/regTable[2][58] , \vrf/regTable[2][59] , \vrf/regTable[2][60] ,
         \vrf/regTable[2][61] , \vrf/regTable[2][62] , \vrf/regTable[2][63] ,
         \vrf/regTable[2][64] , \vrf/regTable[2][65] , \vrf/regTable[2][66] ,
         \vrf/regTable[2][67] , \vrf/regTable[2][68] , \vrf/regTable[2][69] ,
         \vrf/regTable[2][70] , \vrf/regTable[2][71] , \vrf/regTable[2][72] ,
         \vrf/regTable[2][73] , \vrf/regTable[2][74] , \vrf/regTable[2][75] ,
         \vrf/regTable[2][76] , \vrf/regTable[2][77] , \vrf/regTable[2][78] ,
         \vrf/regTable[2][79] , \vrf/regTable[2][80] , \vrf/regTable[2][81] ,
         \vrf/regTable[2][82] , \vrf/regTable[2][83] , \vrf/regTable[2][84] ,
         \vrf/regTable[2][85] , \vrf/regTable[2][86] , \vrf/regTable[2][87] ,
         \vrf/regTable[2][88] , \vrf/regTable[2][89] , \vrf/regTable[2][90] ,
         \vrf/regTable[2][91] , \vrf/regTable[2][92] , \vrf/regTable[2][93] ,
         \vrf/regTable[2][94] , \vrf/regTable[2][95] , \vrf/regTable[2][96] ,
         \vrf/regTable[2][97] , \vrf/regTable[2][98] , \vrf/regTable[2][99] ,
         \vrf/regTable[2][100] , \vrf/regTable[2][101] ,
         \vrf/regTable[2][102] , \vrf/regTable[2][103] ,
         \vrf/regTable[2][104] , \vrf/regTable[2][105] ,
         \vrf/regTable[2][106] , \vrf/regTable[2][107] ,
         \vrf/regTable[2][108] , \vrf/regTable[2][109] ,
         \vrf/regTable[2][110] , \vrf/regTable[2][111] ,
         \vrf/regTable[2][112] , \vrf/regTable[2][113] ,
         \vrf/regTable[2][114] , \vrf/regTable[2][115] ,
         \vrf/regTable[2][116] , \vrf/regTable[2][117] ,
         \vrf/regTable[2][118] , \vrf/regTable[2][119] ,
         \vrf/regTable[2][120] , \vrf/regTable[2][121] ,
         \vrf/regTable[2][122] , \vrf/regTable[2][123] ,
         \vrf/regTable[2][124] , \vrf/regTable[2][125] ,
         \vrf/regTable[2][126] , \vrf/regTable[2][127] ,
         \vrf/regTable[2][128] , \vrf/regTable[2][129] ,
         \vrf/regTable[2][130] , \vrf/regTable[2][131] ,
         \vrf/regTable[2][132] , \vrf/regTable[2][133] ,
         \vrf/regTable[2][134] , \vrf/regTable[2][135] ,
         \vrf/regTable[2][136] , \vrf/regTable[2][137] ,
         \vrf/regTable[2][138] , \vrf/regTable[2][139] ,
         \vrf/regTable[2][140] , \vrf/regTable[2][141] ,
         \vrf/regTable[2][142] , \vrf/regTable[2][143] ,
         \vrf/regTable[2][144] , \vrf/regTable[2][145] ,
         \vrf/regTable[2][146] , \vrf/regTable[2][147] ,
         \vrf/regTable[2][148] , \vrf/regTable[2][149] ,
         \vrf/regTable[2][150] , \vrf/regTable[2][151] ,
         \vrf/regTable[2][152] , \vrf/regTable[2][153] ,
         \vrf/regTable[2][154] , \vrf/regTable[2][155] ,
         \vrf/regTable[2][156] , \vrf/regTable[2][157] ,
         \vrf/regTable[2][158] , \vrf/regTable[2][159] ,
         \vrf/regTable[2][160] , \vrf/regTable[2][161] ,
         \vrf/regTable[2][162] , \vrf/regTable[2][163] ,
         \vrf/regTable[2][164] , \vrf/regTable[2][165] ,
         \vrf/regTable[2][166] , \vrf/regTable[2][167] ,
         \vrf/regTable[2][168] , \vrf/regTable[2][169] ,
         \vrf/regTable[2][170] , \vrf/regTable[2][171] ,
         \vrf/regTable[2][172] , \vrf/regTable[2][173] ,
         \vrf/regTable[2][174] , \vrf/regTable[2][175] ,
         \vrf/regTable[2][176] , \vrf/regTable[2][177] ,
         \vrf/regTable[2][178] , \vrf/regTable[2][179] ,
         \vrf/regTable[2][180] , \vrf/regTable[2][181] ,
         \vrf/regTable[2][182] , \vrf/regTable[2][183] ,
         \vrf/regTable[2][184] , \vrf/regTable[2][185] ,
         \vrf/regTable[2][186] , \vrf/regTable[2][187] ,
         \vrf/regTable[2][188] , \vrf/regTable[2][189] ,
         \vrf/regTable[2][190] , \vrf/regTable[2][191] ,
         \vrf/regTable[2][192] , \vrf/regTable[2][193] ,
         \vrf/regTable[2][194] , \vrf/regTable[2][195] ,
         \vrf/regTable[2][196] , \vrf/regTable[2][197] ,
         \vrf/regTable[2][198] , \vrf/regTable[2][199] ,
         \vrf/regTable[2][200] , \vrf/regTable[2][201] ,
         \vrf/regTable[2][202] , \vrf/regTable[2][203] ,
         \vrf/regTable[2][204] , \vrf/regTable[2][205] ,
         \vrf/regTable[2][206] , \vrf/regTable[2][207] ,
         \vrf/regTable[2][208] , \vrf/regTable[2][209] ,
         \vrf/regTable[2][210] , \vrf/regTable[2][211] ,
         \vrf/regTable[2][212] , \vrf/regTable[2][213] ,
         \vrf/regTable[2][214] , \vrf/regTable[2][215] ,
         \vrf/regTable[2][216] , \vrf/regTable[2][217] ,
         \vrf/regTable[2][218] , \vrf/regTable[2][219] ,
         \vrf/regTable[2][220] , \vrf/regTable[2][221] ,
         \vrf/regTable[2][222] , \vrf/regTable[2][223] ,
         \vrf/regTable[2][224] , \vrf/regTable[2][225] ,
         \vrf/regTable[2][226] , \vrf/regTable[2][227] ,
         \vrf/regTable[2][228] , \vrf/regTable[2][229] ,
         \vrf/regTable[2][230] , \vrf/regTable[2][231] ,
         \vrf/regTable[2][232] , \vrf/regTable[2][233] ,
         \vrf/regTable[2][234] , \vrf/regTable[2][235] ,
         \vrf/regTable[2][236] , \vrf/regTable[2][237] ,
         \vrf/regTable[2][238] , \vrf/regTable[2][239] ,
         \vrf/regTable[2][240] , \vrf/regTable[2][241] ,
         \vrf/regTable[2][242] , \vrf/regTable[2][243] ,
         \vrf/regTable[2][244] , \vrf/regTable[2][245] ,
         \vrf/regTable[2][246] , \vrf/regTable[2][247] ,
         \vrf/regTable[2][248] , \vrf/regTable[2][249] ,
         \vrf/regTable[2][250] , \vrf/regTable[2][251] ,
         \vrf/regTable[2][252] , \vrf/regTable[2][253] ,
         \vrf/regTable[2][254] , \vrf/regTable[2][255] , \vrf/regTable[1][0] ,
         \vrf/regTable[1][1] , \vrf/regTable[1][2] , \vrf/regTable[1][3] ,
         \vrf/regTable[1][4] , \vrf/regTable[1][5] , \vrf/regTable[1][6] ,
         \vrf/regTable[1][7] , \vrf/regTable[1][8] , \vrf/regTable[1][9] ,
         \vrf/regTable[1][10] , \vrf/regTable[1][11] , \vrf/regTable[1][12] ,
         \vrf/regTable[1][13] , \vrf/regTable[1][14] , \vrf/regTable[1][15] ,
         \vrf/regTable[1][16] , \vrf/regTable[1][17] , \vrf/regTable[1][18] ,
         \vrf/regTable[1][19] , \vrf/regTable[1][20] , \vrf/regTable[1][21] ,
         \vrf/regTable[1][22] , \vrf/regTable[1][23] , \vrf/regTable[1][24] ,
         \vrf/regTable[1][25] , \vrf/regTable[1][26] , \vrf/regTable[1][27] ,
         \vrf/regTable[1][28] , \vrf/regTable[1][29] , \vrf/regTable[1][30] ,
         \vrf/regTable[1][31] , \vrf/regTable[1][32] , \vrf/regTable[1][33] ,
         \vrf/regTable[1][34] , \vrf/regTable[1][35] , \vrf/regTable[1][36] ,
         \vrf/regTable[1][37] , \vrf/regTable[1][38] , \vrf/regTable[1][39] ,
         \vrf/regTable[1][40] , \vrf/regTable[1][41] , \vrf/regTable[1][42] ,
         \vrf/regTable[1][43] , \vrf/regTable[1][44] , \vrf/regTable[1][45] ,
         \vrf/regTable[1][46] , \vrf/regTable[1][47] , \vrf/regTable[1][48] ,
         \vrf/regTable[1][49] , \vrf/regTable[1][50] , \vrf/regTable[1][51] ,
         \vrf/regTable[1][52] , \vrf/regTable[1][53] , \vrf/regTable[1][54] ,
         \vrf/regTable[1][55] , \vrf/regTable[1][56] , \vrf/regTable[1][57] ,
         \vrf/regTable[1][58] , \vrf/regTable[1][59] , \vrf/regTable[1][60] ,
         \vrf/regTable[1][61] , \vrf/regTable[1][62] , \vrf/regTable[1][63] ,
         \vrf/regTable[1][64] , \vrf/regTable[1][65] , \vrf/regTable[1][66] ,
         \vrf/regTable[1][67] , \vrf/regTable[1][68] , \vrf/regTable[1][69] ,
         \vrf/regTable[1][70] , \vrf/regTable[1][71] , \vrf/regTable[1][72] ,
         \vrf/regTable[1][73] , \vrf/regTable[1][74] , \vrf/regTable[1][75] ,
         \vrf/regTable[1][76] , \vrf/regTable[1][77] , \vrf/regTable[1][78] ,
         \vrf/regTable[1][79] , \vrf/regTable[1][80] , \vrf/regTable[1][81] ,
         \vrf/regTable[1][82] , \vrf/regTable[1][83] , \vrf/regTable[1][84] ,
         \vrf/regTable[1][85] , \vrf/regTable[1][86] , \vrf/regTable[1][87] ,
         \vrf/regTable[1][88] , \vrf/regTable[1][89] , \vrf/regTable[1][90] ,
         \vrf/regTable[1][91] , \vrf/regTable[1][92] , \vrf/regTable[1][93] ,
         \vrf/regTable[1][94] , \vrf/regTable[1][95] , \vrf/regTable[1][96] ,
         \vrf/regTable[1][97] , \vrf/regTable[1][98] , \vrf/regTable[1][99] ,
         \vrf/regTable[1][100] , \vrf/regTable[1][101] ,
         \vrf/regTable[1][102] , \vrf/regTable[1][103] ,
         \vrf/regTable[1][104] , \vrf/regTable[1][105] ,
         \vrf/regTable[1][106] , \vrf/regTable[1][107] ,
         \vrf/regTable[1][108] , \vrf/regTable[1][109] ,
         \vrf/regTable[1][110] , \vrf/regTable[1][111] ,
         \vrf/regTable[1][112] , \vrf/regTable[1][113] ,
         \vrf/regTable[1][114] , \vrf/regTable[1][115] ,
         \vrf/regTable[1][116] , \vrf/regTable[1][117] ,
         \vrf/regTable[1][118] , \vrf/regTable[1][119] ,
         \vrf/regTable[1][120] , \vrf/regTable[1][121] ,
         \vrf/regTable[1][122] , \vrf/regTable[1][123] ,
         \vrf/regTable[1][124] , \vrf/regTable[1][125] ,
         \vrf/regTable[1][126] , \vrf/regTable[1][127] ,
         \vrf/regTable[1][128] , \vrf/regTable[1][129] ,
         \vrf/regTable[1][130] , \vrf/regTable[1][131] ,
         \vrf/regTable[1][132] , \vrf/regTable[1][133] ,
         \vrf/regTable[1][134] , \vrf/regTable[1][135] ,
         \vrf/regTable[1][136] , \vrf/regTable[1][137] ,
         \vrf/regTable[1][138] , \vrf/regTable[1][139] ,
         \vrf/regTable[1][140] , \vrf/regTable[1][141] ,
         \vrf/regTable[1][142] , \vrf/regTable[1][143] ,
         \vrf/regTable[1][144] , \vrf/regTable[1][145] ,
         \vrf/regTable[1][146] , \vrf/regTable[1][147] ,
         \vrf/regTable[1][148] , \vrf/regTable[1][149] ,
         \vrf/regTable[1][150] , \vrf/regTable[1][151] ,
         \vrf/regTable[1][152] , \vrf/regTable[1][153] ,
         \vrf/regTable[1][154] , \vrf/regTable[1][155] ,
         \vrf/regTable[1][156] , \vrf/regTable[1][157] ,
         \vrf/regTable[1][158] , \vrf/regTable[1][159] ,
         \vrf/regTable[1][160] , \vrf/regTable[1][161] ,
         \vrf/regTable[1][162] , \vrf/regTable[1][163] ,
         \vrf/regTable[1][164] , \vrf/regTable[1][165] ,
         \vrf/regTable[1][166] , \vrf/regTable[1][167] ,
         \vrf/regTable[1][168] , \vrf/regTable[1][169] ,
         \vrf/regTable[1][170] , \vrf/regTable[1][171] ,
         \vrf/regTable[1][172] , \vrf/regTable[1][173] ,
         \vrf/regTable[1][174] , \vrf/regTable[1][175] ,
         \vrf/regTable[1][176] , \vrf/regTable[1][177] ,
         \vrf/regTable[1][178] , \vrf/regTable[1][179] ,
         \vrf/regTable[1][180] , \vrf/regTable[1][181] ,
         \vrf/regTable[1][182] , \vrf/regTable[1][183] ,
         \vrf/regTable[1][184] , \vrf/regTable[1][185] ,
         \vrf/regTable[1][186] , \vrf/regTable[1][187] ,
         \vrf/regTable[1][188] , \vrf/regTable[1][189] ,
         \vrf/regTable[1][190] , \vrf/regTable[1][191] ,
         \vrf/regTable[1][192] , \vrf/regTable[1][193] ,
         \vrf/regTable[1][194] , \vrf/regTable[1][195] ,
         \vrf/regTable[1][196] , \vrf/regTable[1][197] ,
         \vrf/regTable[1][198] , \vrf/regTable[1][199] ,
         \vrf/regTable[1][200] , \vrf/regTable[1][201] ,
         \vrf/regTable[1][202] , \vrf/regTable[1][203] ,
         \vrf/regTable[1][204] , \vrf/regTable[1][205] ,
         \vrf/regTable[1][206] , \vrf/regTable[1][207] ,
         \vrf/regTable[1][208] , \vrf/regTable[1][209] ,
         \vrf/regTable[1][210] , \vrf/regTable[1][211] ,
         \vrf/regTable[1][212] , \vrf/regTable[1][213] ,
         \vrf/regTable[1][214] , \vrf/regTable[1][215] ,
         \vrf/regTable[1][216] , \vrf/regTable[1][217] ,
         \vrf/regTable[1][218] , \vrf/regTable[1][219] ,
         \vrf/regTable[1][220] , \vrf/regTable[1][221] ,
         \vrf/regTable[1][222] , \vrf/regTable[1][223] ,
         \vrf/regTable[1][224] , \vrf/regTable[1][225] ,
         \vrf/regTable[1][226] , \vrf/regTable[1][227] ,
         \vrf/regTable[1][228] , \vrf/regTable[1][229] ,
         \vrf/regTable[1][230] , \vrf/regTable[1][231] ,
         \vrf/regTable[1][232] , \vrf/regTable[1][233] ,
         \vrf/regTable[1][234] , \vrf/regTable[1][235] ,
         \vrf/regTable[1][236] , \vrf/regTable[1][237] ,
         \vrf/regTable[1][238] , \vrf/regTable[1][239] ,
         \vrf/regTable[1][240] , \vrf/regTable[1][241] ,
         \vrf/regTable[1][242] , \vrf/regTable[1][243] ,
         \vrf/regTable[1][244] , \vrf/regTable[1][245] ,
         \vrf/regTable[1][246] , \vrf/regTable[1][247] ,
         \vrf/regTable[1][248] , \vrf/regTable[1][249] ,
         \vrf/regTable[1][250] , \vrf/regTable[1][251] ,
         \vrf/regTable[1][252] , \vrf/regTable[1][253] ,
         \vrf/regTable[1][254] , \vrf/regTable[1][255] , \vrf/regTable[0][0] ,
         \vrf/regTable[0][1] , \vrf/regTable[0][2] , \vrf/regTable[0][3] ,
         \vrf/regTable[0][4] , \vrf/regTable[0][5] , \vrf/regTable[0][6] ,
         \vrf/regTable[0][7] , \vrf/regTable[0][8] , \vrf/regTable[0][9] ,
         \vrf/regTable[0][10] , \vrf/regTable[0][11] , \vrf/regTable[0][12] ,
         \vrf/regTable[0][13] , \vrf/regTable[0][14] , \vrf/regTable[0][15] ,
         \vrf/regTable[0][16] , \vrf/regTable[0][17] , \vrf/regTable[0][18] ,
         \vrf/regTable[0][19] , \vrf/regTable[0][20] , \vrf/regTable[0][21] ,
         \vrf/regTable[0][22] , \vrf/regTable[0][23] , \vrf/regTable[0][24] ,
         \vrf/regTable[0][25] , \vrf/regTable[0][26] , \vrf/regTable[0][27] ,
         \vrf/regTable[0][28] , \vrf/regTable[0][29] , \vrf/regTable[0][30] ,
         \vrf/regTable[0][31] , \vrf/regTable[0][32] , \vrf/regTable[0][33] ,
         \vrf/regTable[0][34] , \vrf/regTable[0][35] , \vrf/regTable[0][36] ,
         \vrf/regTable[0][37] , \vrf/regTable[0][38] , \vrf/regTable[0][39] ,
         \vrf/regTable[0][40] , \vrf/regTable[0][41] , \vrf/regTable[0][42] ,
         \vrf/regTable[0][43] , \vrf/regTable[0][44] , \vrf/regTable[0][45] ,
         \vrf/regTable[0][46] , \vrf/regTable[0][47] , \vrf/regTable[0][48] ,
         \vrf/regTable[0][49] , \vrf/regTable[0][50] , \vrf/regTable[0][51] ,
         \vrf/regTable[0][52] , \vrf/regTable[0][53] , \vrf/regTable[0][54] ,
         \vrf/regTable[0][55] , \vrf/regTable[0][56] , \vrf/regTable[0][57] ,
         \vrf/regTable[0][58] , \vrf/regTable[0][59] , \vrf/regTable[0][60] ,
         \vrf/regTable[0][61] , \vrf/regTable[0][62] , \vrf/regTable[0][63] ,
         \vrf/regTable[0][64] , \vrf/regTable[0][65] , \vrf/regTable[0][66] ,
         \vrf/regTable[0][67] , \vrf/regTable[0][68] , \vrf/regTable[0][69] ,
         \vrf/regTable[0][70] , \vrf/regTable[0][71] , \vrf/regTable[0][72] ,
         \vrf/regTable[0][73] , \vrf/regTable[0][74] , \vrf/regTable[0][75] ,
         \vrf/regTable[0][76] , \vrf/regTable[0][77] , \vrf/regTable[0][78] ,
         \vrf/regTable[0][79] , \vrf/regTable[0][80] , \vrf/regTable[0][81] ,
         \vrf/regTable[0][82] , \vrf/regTable[0][83] , \vrf/regTable[0][84] ,
         \vrf/regTable[0][85] , \vrf/regTable[0][86] , \vrf/regTable[0][87] ,
         \vrf/regTable[0][88] , \vrf/regTable[0][89] , \vrf/regTable[0][90] ,
         \vrf/regTable[0][91] , \vrf/regTable[0][92] , \vrf/regTable[0][93] ,
         \vrf/regTable[0][94] , \vrf/regTable[0][95] , \vrf/regTable[0][96] ,
         \vrf/regTable[0][97] , \vrf/regTable[0][98] , \vrf/regTable[0][99] ,
         \vrf/regTable[0][100] , \vrf/regTable[0][101] ,
         \vrf/regTable[0][102] , \vrf/regTable[0][103] ,
         \vrf/regTable[0][104] , \vrf/regTable[0][105] ,
         \vrf/regTable[0][106] , \vrf/regTable[0][107] ,
         \vrf/regTable[0][108] , \vrf/regTable[0][109] ,
         \vrf/regTable[0][110] , \vrf/regTable[0][111] ,
         \vrf/regTable[0][112] , \vrf/regTable[0][113] ,
         \vrf/regTable[0][114] , \vrf/regTable[0][115] ,
         \vrf/regTable[0][116] , \vrf/regTable[0][117] ,
         \vrf/regTable[0][118] , \vrf/regTable[0][119] ,
         \vrf/regTable[0][120] , \vrf/regTable[0][121] ,
         \vrf/regTable[0][122] , \vrf/regTable[0][123] ,
         \vrf/regTable[0][124] , \vrf/regTable[0][125] ,
         \vrf/regTable[0][126] , \vrf/regTable[0][127] ,
         \vrf/regTable[0][128] , \vrf/regTable[0][129] ,
         \vrf/regTable[0][130] , \vrf/regTable[0][131] ,
         \vrf/regTable[0][132] , \vrf/regTable[0][133] ,
         \vrf/regTable[0][134] , \vrf/regTable[0][135] ,
         \vrf/regTable[0][136] , \vrf/regTable[0][137] ,
         \vrf/regTable[0][138] , \vrf/regTable[0][139] ,
         \vrf/regTable[0][140] , \vrf/regTable[0][141] ,
         \vrf/regTable[0][142] , \vrf/regTable[0][143] ,
         \vrf/regTable[0][144] , \vrf/regTable[0][145] ,
         \vrf/regTable[0][146] , \vrf/regTable[0][147] ,
         \vrf/regTable[0][148] , \vrf/regTable[0][149] ,
         \vrf/regTable[0][150] , \vrf/regTable[0][151] ,
         \vrf/regTable[0][152] , \vrf/regTable[0][153] ,
         \vrf/regTable[0][154] , \vrf/regTable[0][155] ,
         \vrf/regTable[0][156] , \vrf/regTable[0][157] ,
         \vrf/regTable[0][158] , \vrf/regTable[0][159] ,
         \vrf/regTable[0][160] , \vrf/regTable[0][161] ,
         \vrf/regTable[0][162] , \vrf/regTable[0][163] ,
         \vrf/regTable[0][164] , \vrf/regTable[0][165] ,
         \vrf/regTable[0][166] , \vrf/regTable[0][167] ,
         \vrf/regTable[0][168] , \vrf/regTable[0][169] ,
         \vrf/regTable[0][170] , \vrf/regTable[0][171] ,
         \vrf/regTable[0][172] , \vrf/regTable[0][173] ,
         \vrf/regTable[0][174] , \vrf/regTable[0][175] ,
         \vrf/regTable[0][176] , \vrf/regTable[0][177] ,
         \vrf/regTable[0][178] , \vrf/regTable[0][179] ,
         \vrf/regTable[0][180] , \vrf/regTable[0][181] ,
         \vrf/regTable[0][182] , \vrf/regTable[0][183] ,
         \vrf/regTable[0][184] , \vrf/regTable[0][185] ,
         \vrf/regTable[0][186] , \vrf/regTable[0][187] ,
         \vrf/regTable[0][188] , \vrf/regTable[0][189] ,
         \vrf/regTable[0][190] , \vrf/regTable[0][191] ,
         \vrf/regTable[0][192] , \vrf/regTable[0][193] ,
         \vrf/regTable[0][194] , \vrf/regTable[0][195] ,
         \vrf/regTable[0][196] , \vrf/regTable[0][197] ,
         \vrf/regTable[0][198] , \vrf/regTable[0][199] ,
         \vrf/regTable[0][200] , \vrf/regTable[0][201] ,
         \vrf/regTable[0][202] , \vrf/regTable[0][203] ,
         \vrf/regTable[0][204] , \vrf/regTable[0][205] ,
         \vrf/regTable[0][206] , \vrf/regTable[0][207] ,
         \vrf/regTable[0][208] , \vrf/regTable[0][209] ,
         \vrf/regTable[0][210] , \vrf/regTable[0][211] ,
         \vrf/regTable[0][212] , \vrf/regTable[0][213] ,
         \vrf/regTable[0][214] , \vrf/regTable[0][215] ,
         \vrf/regTable[0][216] , \vrf/regTable[0][217] ,
         \vrf/regTable[0][218] , \vrf/regTable[0][219] ,
         \vrf/regTable[0][220] , \vrf/regTable[0][221] ,
         \vrf/regTable[0][222] , \vrf/regTable[0][223] ,
         \vrf/regTable[0][224] , \vrf/regTable[0][225] ,
         \vrf/regTable[0][226] , \vrf/regTable[0][227] ,
         \vrf/regTable[0][228] , \vrf/regTable[0][229] ,
         \vrf/regTable[0][230] , \vrf/regTable[0][231] ,
         \vrf/regTable[0][232] , \vrf/regTable[0][233] ,
         \vrf/regTable[0][234] , \vrf/regTable[0][235] ,
         \vrf/regTable[0][236] , \vrf/regTable[0][237] ,
         \vrf/regTable[0][238] , \vrf/regTable[0][239] ,
         \vrf/regTable[0][240] , \vrf/regTable[0][241] ,
         \vrf/regTable[0][242] , \vrf/regTable[0][243] ,
         \vrf/regTable[0][244] , \vrf/regTable[0][245] ,
         \vrf/regTable[0][246] , \vrf/regTable[0][247] ,
         \vrf/regTable[0][248] , \vrf/regTable[0][249] ,
         \vrf/regTable[0][250] , \vrf/regTable[0][251] ,
         \vrf/regTable[0][252] , \vrf/regTable[0][253] ,
         \vrf/regTable[0][254] , \vrf/regTable[0][255] , \vrf/N14 , \vrf/N13 ,
         \vrf/N12 , \vrf/N11 , \vrf/N10 , \vrf/N9 , \srf/N59 , \srf/N58 ,
         \srf/N57 , \srf/N56 , \srf/N55 , \srf/N54 , \srf/N53 , \srf/N52 ,
         \srf/N51 , \srf/N50 , \srf/N49 , \srf/N48 , \srf/N47 , \srf/N46 ,
         \srf/N45 , \srf/N44 , \srf/N43 , \srf/N42 , \srf/N41 , \srf/N40 ,
         \srf/N39 , \srf/N38 , \srf/N37 , \srf/N36 , \srf/N35 , \srf/N34 ,
         \srf/N33 , \srf/N32 , \srf/N31 , \srf/N30 , \srf/N29 , \srf/N28 ,
         \srf/N27 , \srf/N26 , \srf/N25 , \srf/N24 , \srf/N23 , \srf/N22 ,
         \srf/N21 , \srf/N20 , \srf/regTable[7][0] , \srf/regTable[7][1] ,
         \srf/regTable[7][2] , \srf/regTable[7][3] , \srf/regTable[7][4] ,
         \srf/regTable[7][5] , \srf/regTable[7][6] , \srf/regTable[7][7] ,
         \srf/regTable[7][8] , \srf/regTable[7][9] , \srf/regTable[7][10] ,
         \srf/regTable[7][11] , \srf/regTable[7][12] , \srf/regTable[7][13] ,
         \srf/regTable[7][14] , \srf/regTable[7][15] , \srf/regTable[6][0] ,
         \srf/regTable[6][1] , \srf/regTable[6][2] , \srf/regTable[6][3] ,
         \srf/regTable[6][4] , \srf/regTable[6][5] , \srf/regTable[6][6] ,
         \srf/regTable[6][7] , \srf/regTable[6][8] , \srf/regTable[6][9] ,
         \srf/regTable[6][10] , \srf/regTable[6][11] , \srf/regTable[6][12] ,
         \srf/regTable[6][13] , \srf/regTable[6][14] , \srf/regTable[6][15] ,
         \srf/regTable[5][0] , \srf/regTable[5][1] , \srf/regTable[5][2] ,
         \srf/regTable[5][3] , \srf/regTable[5][4] , \srf/regTable[5][5] ,
         \srf/regTable[5][6] , \srf/regTable[5][7] , \srf/regTable[5][8] ,
         \srf/regTable[5][9] , \srf/regTable[5][10] , \srf/regTable[5][11] ,
         \srf/regTable[5][12] , \srf/regTable[5][13] , \srf/regTable[5][14] ,
         \srf/regTable[5][15] , \srf/regTable[4][0] , \srf/regTable[4][1] ,
         \srf/regTable[4][2] , \srf/regTable[4][3] , \srf/regTable[4][4] ,
         \srf/regTable[4][5] , \srf/regTable[4][6] , \srf/regTable[4][7] ,
         \srf/regTable[4][8] , \srf/regTable[4][9] , \srf/regTable[4][10] ,
         \srf/regTable[4][11] , \srf/regTable[4][12] , \srf/regTable[4][13] ,
         \srf/regTable[4][14] , \srf/regTable[4][15] , \srf/regTable[3][0] ,
         \srf/regTable[3][1] , \srf/regTable[3][2] , \srf/regTable[3][3] ,
         \srf/regTable[3][4] , \srf/regTable[3][5] , \srf/regTable[3][6] ,
         \srf/regTable[3][7] , \srf/regTable[3][8] , \srf/regTable[3][9] ,
         \srf/regTable[3][10] , \srf/regTable[3][11] , \srf/regTable[3][12] ,
         \srf/regTable[3][13] , \srf/regTable[3][14] , \srf/regTable[3][15] ,
         \srf/regTable[2][0] , \srf/regTable[2][1] , \srf/regTable[2][2] ,
         \srf/regTable[2][3] , \srf/regTable[2][4] , \srf/regTable[2][5] ,
         \srf/regTable[2][6] , \srf/regTable[2][7] , \srf/regTable[2][8] ,
         \srf/regTable[2][9] , \srf/regTable[2][10] , \srf/regTable[2][11] ,
         \srf/regTable[2][12] , \srf/regTable[2][13] , \srf/regTable[2][14] ,
         \srf/regTable[2][15] , \srf/regTable[1][0] , \srf/regTable[1][1] ,
         \srf/regTable[1][2] , \srf/regTable[1][3] , \srf/regTable[1][4] ,
         \srf/regTable[1][5] , \srf/regTable[1][6] , \srf/regTable[1][7] ,
         \srf/regTable[1][8] , \srf/regTable[1][9] , \srf/regTable[1][10] ,
         \srf/regTable[1][11] , \srf/regTable[1][12] , \srf/regTable[1][13] ,
         \srf/regTable[1][14] , \srf/regTable[1][15] , \srf/regTable[0][0] ,
         \srf/regTable[0][1] , \srf/regTable[0][2] , \srf/regTable[0][3] ,
         \srf/regTable[0][4] , \srf/regTable[0][5] , \srf/regTable[0][6] ,
         \srf/regTable[0][7] , \srf/regTable[0][8] , \srf/regTable[0][9] ,
         \srf/regTable[0][10] , \srf/regTable[0][11] , \srf/regTable[0][12] ,
         \srf/regTable[0][13] , \srf/regTable[0][14] , \srf/regTable[0][15] ,
         \srf/N17 , \srf/N16 , \srf/N15 , \alu/N1019 , \alu/N1018 ,
         \alu/N1017 , \alu/N1016 , \alu/N1015 , \alu/N1014 , \alu/N1013 ,
         \alu/N1012 , \alu/N1011 , \alu/N1010 , \alu/N1009 , \alu/N1008 ,
         \alu/N1007 , \alu/N1006 , \alu/N1005 , \alu/N1004 , \alu/N999 ,
         \alu/N997 , \alu/N991 , \alu/N990 , \alu/N989 , \alu/N988 ,
         \alu/N987 , \alu/N986 , \alu/N985 , \alu/N984 , \alu/N983 ,
         \alu/N982 , \alu/N851 , \alu/N850 , \alu/N849 , \alu/N848 ,
         \alu/N847 , \alu/N846 , \alu/N845 , \alu/N844 , \alu/N843 ,
         \alu/N842 , \alu/N841 , \alu/N840 , \alu/N839 , \alu/N836 ,
         \alu/N835 , \alu/N834 , \alu/N833 , \alu/N814 , \alu/N665 ,
         \alu/N664 , \alu/N663 , \alu/N662 , \alu/N661 , \alu/N660 ,
         \alu/N659 , \alu/N658 , \alu/N657 , \alu/N656 , \alu/N655 ,
         \alu/N654 , \alu/N653 , \alu/N652 , \alu/N651 , \alu/N634 ,
         \alu/N610 , \alu/N609 , \alu/N608 , \alu/N607 , \alu/N606 ,
         \alu/N605 , \alu/N604 , \alu/N603 , \alu/N602 , \alu/N601 ,
         \alu/N600 , \alu/N579 , \alu/N543 , \alu/N542 , \alu/N541 ,
         \alu/N540 , \alu/N539 , \alu/N529 , \alu/N521 , \alu/N520 ,
         \alu/N519 , \alu/N477 , \alu/N476 , \alu/N475 , \alu/N474 ,
         \alu/N473 , \alu/N472 , \alu/N471 , \alu/N470 , \alu/N469 ,
         \alu/N468 , \alu/N467 , \alu/N466 , \alu/N465 , \alu/N464 ,
         \alu/N456 , \alu/N455 , \alu/N454 , \alu/N453 , \alu/N452 ,
         \alu/N451 , \alu/N450 , \alu/N449 , \alu/N448 , \alu/N447 ,
         \alu/N446 , \alu/N443 , \alu/N442 , \alu/N441 , \alu/N440 ,
         \alu/N439 , \alu/N438 , \alu/N433 , \alu/N432 , \alu/N431 ,
         \alu/N424 , \alu/N423 , \alu/N422 , \alu/N421 , \alu/N420 ,
         \alu/N419 , \alu/N418 , \alu/N417 , \alu/N416 , \alu/N415 ,
         \alu/N414 , \alu/N413 , \alu/N412 , \alu/N411 , \alu/N410 ,
         \alu/N409 , \alu/N408 , \alu/N407 , \alu/N406 , \alu/N385 ,
         \alu/N376 , \alu/N338 , \alu/N337 , \alu/N336 , \alu/N335 ,
         \alu/N334 , \alu/N333 , \alu/N332 , \alu/N331 , \alu/N330 ,
         \alu/N329 , \alu/N328 , \alu/N327 , \alu/N326 , \alu/N312 ,
         \alu/N311 , \alu/N310 , \alu/N309 , \alu/N308 , \alu/N307 ,
         \alu/N293 , \alu/N292 , \alu/N291 , \alu/N290 , \alu/N289 ,
         \alu/N288 , \alu/N287 , \alu/N286 , \alu/N285 , \alu/N284 ,
         \alu/N283 , \alu/N282 , \alu/N281 , \alu/N226 , \alu/N225 ,
         \alu/N224 , \alu/N223 , \alu/N222 , \alu/N221 , \alu/N220 ,
         \alu/N219 , \alu/N218 , \alu/N217 , \alu/N216 , \alu/N215 ,
         \alu/N214 , \alu/N213 , \alu/N212 , \alu/N211 , \alu/N210 ,
         \alu/N209 , \alu/N208 , \alu/N207 , \alu/N206 , \alu/N205 ,
         \alu/N204 , \alu/N203 , \alu/N202 , \alu/N201 , \alu/N117 ,
         \alu/N116 , \alu/N115 , \alu/N114 , \alu/N113 , \alu/N112 ,
         \alu/N111 , \alu/N110 , \alu/N109 , \alu/N108 , \alu/N107 ,
         \alu/N106 , \alu/N105 , \alu/N104 , \alu/N103 , \alu/N102 ,
         \alu/N101 , \alu/N100 , \alu/N99 , \alu/N98 , \alu/N97 , \alu/N96 ,
         \alu/N95 , \alu/N94 , \alu/N93 , \alu/N92 , \alu/N88 , \alu/N87 ,
         \*Logic0* , \alu/*Logic1* , n214, n215, n216, n217, n218, n219,
         \U3/U6/Z_15 , \U3/U6/Z_16 , \U3/U6/Z_17 , \U3/U6/Z_18 , \U3/U6/Z_19 ,
         \U3/U6/Z_20 , \U3/U6/Z_21 , \U3/U6/Z_22 , \U3/U6/Z_23 , \U3/U6/Z_24 ,
         \U3/U6/Z_25 , \U3/U7/Z_0 , \U3/U7/Z_1 , \U3/U7/Z_2 , \U3/U7/Z_3 ,
         \U3/U7/Z_4 , \U3/U7/Z_5 , \U3/U7/Z_6 , \U3/U7/Z_7 , \U3/U7/Z_8 ,
         \U3/U7/Z_9 , \U3/U7/Z_10 , \U3/U7/Z_11 , \U3/U7/Z_12 , \U3/U7/Z_13 ,
         \U3/U7/Z_14 , \U3/U7/Z_15 , \U3/U7/Z_16 , \U3/U7/Z_17 , \U3/U7/Z_18 ,
         \U3/U7/Z_19 , \U3/U7/Z_20 , \U3/U7/Z_21 , \U3/U7/Z_22 , \U3/U7/Z_23 ,
         \U3/U7/Z_24 , \U3/U7/Z_25 , \U3/U8/Z_0 , \U3/U13/Z_0 , \U3/U13/Z_1 ,
         \U3/U13/Z_2 , \U3/U13/Z_3 , \U3/U13/Z_4 , \U3/U13/Z_5 , \U3/U13/Z_6 ,
         \U3/U13/Z_7 , \U3/U13/Z_8 , \U3/U13/Z_9 , \U3/U13/Z_10 ,
         \U3/U13/Z_11 , \U3/U13/Z_12 , \U3/U13/Z_13 , \U3/U13/Z_14 ,
         \U3/U13/Z_15 , \U3/U14/Z_0 , \U3/U14/Z_1 , \U3/U14/Z_2 , \U3/U14/Z_3 ,
         \U3/U14/Z_4 , \U3/U16/Z_0 , \U3/U16/Z_1 , \U3/U16/Z_2 , \U3/U16/Z_3 ,
         \U3/U16/Z_4 , \U3/U17/Z_0 , \U3/U17/Z_1 , \U3/U17/Z_2 , \U3/U17/Z_3 ,
         \U3/U19/Z_0 , \U3/U19/Z_1 , \U3/U19/Z_2 , \U3/U19/Z_3 , \U3/U22/Z_0 ,
         \U3/U22/Z_1 , \U3/U22/Z_2 , \U3/U22/Z_3 , \U3/U22/Z_4 , \U3/U22/Z_5 ,
         \U3/U23/Z_0 , \U3/U23/Z_1 , \U3/U23/Z_2 , \U3/U23/Z_3 , \U3/U24/Z_0 ,
         \U3/U25/Z_15 , \U3/U25/Z_16 , \U3/U25/Z_17 , \U3/U25/Z_18 ,
         \U3/U25/Z_19 , \U3/U25/Z_20 , \U3/U25/Z_21 , \U3/U25/Z_22 ,
         \U3/U25/Z_23 , \U3/U25/Z_24 , \U3/U25/Z_25 , \U3/U26/Z_0 ,
         \U3/U26/Z_1 , \U3/U26/Z_2 , \U3/U26/Z_3 , \U3/U26/Z_4 , \U3/U26/Z_5 ,
         \U3/U26/Z_6 , \U3/U26/Z_7 , \U3/U26/Z_8 , \U3/U26/Z_9 , \U3/U26/Z_10 ,
         \U3/U26/Z_11 , \U3/U26/Z_12 , \U3/U26/Z_13 , \U3/U26/Z_14 ,
         \U3/U26/Z_15 , \U3/U26/Z_16 , \U3/U26/Z_17 , \U3/U26/Z_18 ,
         \U3/U26/Z_19 , \U3/U26/Z_20 , \U3/U26/Z_21 , \U3/U26/Z_22 ,
         \U3/U26/Z_23 , \U3/U26/Z_24 , \U3/U26/Z_25 , \U3/U27/Z_0 ,
         \U3/U29/Z_0 , \U3/U29/Z_1 , \U3/U29/Z_2 , \U3/U29/Z_3 , \U3/U29/Z_4 ,
         \U3/U30/Z_0 , \U3/U30/Z_1 , \U3/U30/Z_2 , \U3/U30/Z_3 , \U3/U30/Z_4 ,
         \U3/U31/Z_0 , \U3/U32/Z_0 , n1461, n2522, n3262, n3266, n3368, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476;
  wire   [255:0] vectorData1;
  wire   [255:0] vectorData2;
  wire   [15:0] scalarWrData;
  wire   [15:0] scalarData1;
  wire   [15:0] scalarData2;
  wire   [255:0] op1;
  wire   [255:0] op2;
  wire   [3:0] func;
  wire   [255:0] result;
  wire   [15:0] instrIn;
  wire   [2:0] addrDst;
  wire   [3:0] code;
  wire   [3:0] state;
  wire   [4:0] cycles;
  wire   [15:0] scalarToLoad;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90;

  LHQD4BWP \cycles_reg[4]  ( .E(N4064), .D(N4069), .Q(cycles[4]) );
  LHQD4BWP \cycles_reg[3]  ( .E(N4064), .D(N4068), .Q(cycles[3]) );
  LHQD4BWP \cycles_reg[0]  ( .E(N4064), .D(N4065), .Q(cycles[0]) );
  LHQD4BWP \cycles_reg[1]  ( .E(N4064), .D(N4066), .Q(cycles[1]) );
  LHQD4BWP \cycles_reg[2]  ( .E(N4064), .D(N4067), .Q(cycles[2]) );
  CVP14_DW01_addsub_0 r1183 ( .A({\U3/U16/Z_4 , \U3/U16/Z_3 , \U3/U16/Z_2 , 
        \U3/U16/Z_1 , \U3/U16/Z_0 }), .B({\*Logic0* , \U3/U17/Z_3 , 
        \U3/U17/Z_2 , \U3/U17/Z_1 , \U3/U17/Z_0 }), .CI(\*Logic0* ), .ADD_SUB(
        n7440), .SUM({N3436, N3435, N3434, N3433, N3432}) );
  CVP14_DW01_ash_0 sll_485_C216 ( .A({n7449, N1610, n7448, n7447, n7446, n7445, 
        n7444, n7443, n7442, N1602, N1601, N1600}), .DATA_TC(\*Logic0* ), .SH(
        {n7439, N1660, n7441, N1681}), .SH_TC(\*Logic0* ), .B({N1691, N1690, 
        N1689, N1688, N1687, N1686, N1685, N1684, N1683, N1682, 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1}) );
  CVP14_DW01_decode_0 r806 ( .A(cycles), .B({SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, N1108, N1107, 
        N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, 
        N1096, N1095, N1094}) );
  CVP14_DW01_ash_1 r803 ( .A({\*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , n7476, result[15:0]}), .DATA_TC(\*Logic0* ), .SH({cycles, 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* }), .SH_TC(\*Logic0* ), 
        .B({N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, 
        N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, 
        N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, 
        N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, 
        N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, 
        N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, 
        N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, 
        N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, 
        N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, 
        N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, 
        N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, 
        N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, 
        N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, 
        N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, 
        N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, 
        N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, 
        N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, 
        N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, 
        N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, 
        N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, 
        N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, 
        N321, N320, N319, N318, N317}) );
  CVP14_DW01_decode_1 r801 ( .A(cycles), .B({SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, N267, N266, N265, 
        N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253}) );
  CVP14_DW01_ash_2 sll_264 ( .A({\*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , DataIn}), .DATA_TC(\*Logic0* ), 
        .SH({N2626, N2626, N2626, N2626, N2626, N2626, N2626, N2626, N2626, 
        N2626, N2626, N2626, N2626, N2626, N2626, N2626, N2626, N2626, N2626, 
        N2626, N2626, N2626, N2626, N1565, N1564, N1563, N1562, N1561, 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* }), .SH_TC(\*Logic0* ), 
        .B({N2882, N2881, N2880, N2879, N2878, N2877, N2876, N2875, N2874, 
        N2873, N2872, N2871, N2870, N2869, N2868, N2867, N2866, N2865, N2864, 
        N2863, N2862, N2861, N2860, N2859, N2858, N2857, N2856, N2855, N2854, 
        N2853, N2852, N2851, N2850, N2849, N2848, N2847, N2846, N2845, N2844, 
        N2843, N2842, N2841, N2840, N2839, N2838, N2837, N2836, N2835, N2834, 
        N2833, N2832, N2831, N2830, N2829, N2828, N2827, N2826, N2825, N2824, 
        N2823, N2822, N2821, N2820, N2819, N2818, N2817, N2816, N2815, N2814, 
        N2813, N2812, N2811, N2810, N2809, N2808, N2807, N2806, N2805, N2804, 
        N2803, N2802, N2801, N2800, N2799, N2798, N2797, N2796, N2795, N2794, 
        N2793, N2792, N2791, N2790, N2789, N2788, N2787, N2786, N2785, N2784, 
        N2783, N2782, N2781, N2780, N2779, N2778, N2777, N2776, N2775, N2774, 
        N2773, N2772, N2771, N2770, N2769, N2768, N2767, N2766, N2765, N2764, 
        N2763, N2762, N2761, N2760, N2759, N2758, N2757, N2756, N2755, N2754, 
        N2753, N2752, N2751, N2750, N2749, N2748, N2747, N2746, N2745, N2744, 
        N2743, N2742, N2741, N2740, N2739, N2738, N2737, N2736, N2735, N2734, 
        N2733, N2732, N2731, N2730, N2729, N2728, N2727, N2726, N2725, N2724, 
        N2723, N2722, N2721, N2720, N2719, N2718, N2717, N2716, N2715, N2714, 
        N2713, N2712, N2711, N2710, N2709, N2708, N2707, N2706, N2705, N2704, 
        N2703, N2702, N2701, N2700, N2699, N2698, N2697, N2696, N2695, N2694, 
        N2693, N2692, N2691, N2690, N2689, N2688, N2687, N2686, N2685, N2684, 
        N2683, N2682, N2681, N2680, N2679, N2678, N2677, N2676, N2675, N2674, 
        N2673, N2672, N2671, N2670, N2669, N2668, N2667, N2666, N2665, N2664, 
        N2663, N2662, N2661, N2660, N2659, N2658, N2657, N2656, N2655, N2654, 
        N2653, N2652, N2651, N2650, N2649, N2648, N2647, N2646, N2645, N2644, 
        N2643, N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635, N2634, 
        N2633, N2632, N2631, N2630, N2629, N2628, N2627}) );
  CVP14_DW01_inc_1 add_461_C216 ( .A({\*Logic0* , N1537, N1536, N1535, N1534, 
        N1533, N1532, N1531, N1530, N1529, N1528, N1527, n7455, n7454, N1524, 
        N1523, N1522, N1521, N1520, N1519, n7453, n7452, n7451, n7450, N1514, 
        N1513, N1512}), .SUM({N1558, N1557, N1556, N1555, N1554, N1553, N1552, 
        N1551, N1550, N1549, N1548, N1547, N1546, N1545, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48}) );
  CVP14_DW01_ash_3 sll_450_C216 ( .A({N1419, N1418, N1417, N1416, N1415, N1414, 
        N1413, N1412, N1411, N1410, N1409, N1408, N1407}), .DATA_TC(\*Logic0* ), .SH({N1457, N1466, n7457, N1487}), .SH_TC(\*Logic0* ), .B({N1500, N1499, 
        N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, 
        N1488}) );
  CVP14_DW01_addsub_1 r156 ( .A({\U3/U13/Z_15 , \U3/U13/Z_14 , \U3/U13/Z_13 , 
        \U3/U13/Z_12 , \U3/U13/Z_11 , \U3/U13/Z_10 , \U3/U13/Z_9 , 
        \U3/U13/Z_8 , \U3/U13/Z_7 , \U3/U13/Z_6 , \U3/U13/Z_5 , \U3/U13/Z_4 , 
        \U3/U13/Z_3 , \U3/U13/Z_2 , \U3/U13/Z_1 , \U3/U13/Z_0 }), .B({
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \U3/U14/Z_4 , \U3/U14/Z_3 , \U3/U14/Z_2 , \U3/U14/Z_1 , \U3/U14/Z_0 }), 
        .CI(\*Logic0* ), .ADD_SUB(n7456), .SUM({N222, N221, N220, N219, N218, 
        N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207}) );
  CVP14_DW01_addsub_2 r148 ( .A({\*Logic0* , \U3/U6/Z_25 , \U3/U6/Z_24 , 
        \U3/U6/Z_23 , \U3/U6/Z_22 , \U3/U6/Z_21 , \U3/U6/Z_20 , \U3/U6/Z_19 , 
        \U3/U6/Z_18 , \U3/U6/Z_17 , \U3/U6/Z_16 , \U3/U6/Z_15 , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* }), .B({\*Logic0* , \U3/U7/Z_25 , \U3/U7/Z_24 , 
        \U3/U7/Z_23 , \U3/U7/Z_22 , \U3/U7/Z_21 , \U3/U7/Z_20 , \U3/U7/Z_19 , 
        \U3/U7/Z_18 , \U3/U7/Z_17 , \U3/U7/Z_16 , \U3/U7/Z_15 , \U3/U7/Z_14 , 
        \U3/U7/Z_13 , \U3/U7/Z_12 , \U3/U7/Z_11 , \U3/U7/Z_10 , \U3/U7/Z_9 , 
        \U3/U7/Z_8 , \U3/U7/Z_7 , \U3/U7/Z_6 , \U3/U7/Z_5 , \U3/U7/Z_4 , 
        \U3/U7/Z_3 , \U3/U7/Z_2 , \U3/U7/Z_1 , \U3/U7/Z_0 }), .CI(\*Logic0* ), 
        .ADD_SUB(\U3/U8/Z_0 ), .SUM({N1280, N1419, N1418, N1417, N1416, N1415, 
        N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1266, N1265, 
        N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, 
        N1254}) );
  CVP14_DW_rash_0 srl_430_C216 ( .A({N1169, result[9:0], \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* }), .DATA_TC(\*Logic0* ), .SH({N1167, N1166, 
        N1165, N1164, N1163}), .SH_TC(\*Logic0* ), .B({N1307, N1306, N1305, 
        N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, 
        N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, 
        N1284, N1283, N1282}) );
  CVP14_DW_rash_1 srl_424_C216 ( .A({N1168, scalarToLoad[9:0], \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* }), .DATA_TC(\*Logic0* ), .SH({N1167, N1166, 
        N1165, N1164, N1163}), .SH_TC(\*Logic0* ), .B({N1198, N1197, N1196, 
        N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, 
        N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, 
        N1175, N1174, N1173}) );
  CVP14_DW01_ash_4 \alu/sll_191_C23  ( .A({n7460, \alu/N529 , n7467, n7466, 
        n7465, n7464, n7463, n7462, n7461, \alu/N521 , \alu/N520 , \alu/N519 }), .DATA_TC(\*Logic0* ), .SH({n7458, \alu/N579 , n7459, \alu/N600 }), .SH_TC(
        \*Logic0* ), .B({\alu/N610 , \alu/N609 , \alu/N608 , \alu/N607 , 
        \alu/N606 , \alu/N605 , \alu/N604 , \alu/N603 , \alu/N602 , \alu/N601 , 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50}) );
  CVP14_DW01_addsub_3 r1196 ( .A({\U3/U22/Z_5 , \U3/U22/Z_4 , \U3/U22/Z_3 , 
        \U3/U22/Z_2 , \U3/U22/Z_1 , \U3/U22/Z_0 }), .B({\*Logic0* , \*Logic0* , 
        \U3/U23/Z_3 , \U3/U23/Z_2 , \U3/U23/Z_1 , \U3/U23/Z_0 }), .CI(
        \*Logic0* ), .ADD_SUB(\U3/U24/Z_0 ), .SUM({\alu/N997 , \alu/N543 , 
        \alu/N542 , \alu/N541 , \alu/N540 , \alu/N539 }) );
  CVP14_DW01_inc_2 \alu/add_167_C23  ( .A({\*Logic0* , \alu/N456 , \alu/N455 , 
        \alu/N454 , \alu/N453 , \alu/N452 , \alu/N451 , \alu/N450 , \alu/N449 , 
        \alu/N448 , \alu/N447 , \alu/N446 , n7468, n7469, \alu/N443 , 
        \alu/N442 , \alu/N441 , \alu/N440 , \alu/N439 , \alu/N438 , n7473, 
        n7472, n7471, n7470, \alu/N433 , \alu/N432 , \alu/N431 }), .SUM({
        \alu/N477 , \alu/N476 , \alu/N475 , \alu/N474 , \alu/N473 , \alu/N472 , 
        \alu/N471 , \alu/N470 , \alu/N469 , \alu/N468 , \alu/N467 , \alu/N466 , 
        \alu/N465 , \alu/N464 , SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63}) );
  CVP14_DW01_ash_5 \alu/sll_156_C23  ( .A({\alu/N338 , \alu/N337 , \alu/N336 , 
        \alu/N335 , \alu/N334 , \alu/N333 , \alu/N332 , \alu/N331 , \alu/N330 , 
        \alu/N329 , \alu/N328 , \alu/N327 , \alu/N326 }), .DATA_TC(\*Logic0* ), 
        .SH({\alu/N376 , \alu/N385 , n7475, \alu/N406 }), .SH_TC(\*Logic0* ), 
        .B({\alu/N419 , \alu/N418 , \alu/N417 , \alu/N416 , \alu/N415 , 
        \alu/N414 , \alu/N413 , \alu/N412 , \alu/N411 , \alu/N410 , \alu/N409 , 
        \alu/N408 , \alu/N407 }) );
  CVP14_DW01_addsub_5 r1207 ( .A({\alu/N312 , \alu/N311 , \alu/N310 , 
        \alu/N309 , \alu/N308 }), .B({\*Logic0* , \U3/U19/Z_3 , \U3/U19/Z_2 , 
        \U3/U19/Z_1 , \U3/U19/Z_0 }), .CI(\*Logic0* ), .ADD_SUB(n7474), .SUM({
        \alu/N424 , \alu/N423 , \alu/N422 , \alu/N421 , \alu/N420 }) );
  CVP14_DW01_addsub_6 r1208 ( .A({\*Logic0* , \U3/U25/Z_25 , \U3/U25/Z_24 , 
        \U3/U25/Z_23 , \U3/U25/Z_22 , \U3/U25/Z_21 , \U3/U25/Z_20 , 
        \U3/U25/Z_19 , \U3/U25/Z_18 , \U3/U25/Z_17 , \U3/U25/Z_16 , 
        \U3/U25/Z_15 , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* }), .B({
        \*Logic0* , \U3/U26/Z_25 , \U3/U26/Z_24 , \U3/U26/Z_23 , \U3/U26/Z_22 , 
        \U3/U26/Z_21 , \U3/U26/Z_20 , \U3/U26/Z_19 , \U3/U26/Z_18 , 
        \U3/U26/Z_17 , \U3/U26/Z_16 , \U3/U26/Z_15 , \U3/U26/Z_14 , 
        \U3/U26/Z_13 , \U3/U26/Z_12 , \U3/U26/Z_11 , \U3/U26/Z_10 , 
        \U3/U26/Z_9 , \U3/U26/Z_8 , \U3/U26/Z_7 , \U3/U26/Z_6 , \U3/U26/Z_5 , 
        \U3/U26/Z_4 , \U3/U26/Z_3 , \U3/U26/Z_2 , \U3/U26/Z_1 , \U3/U26/Z_0 }), 
        .CI(\*Logic0* ), .ADD_SUB(\U3/U27/Z_0 ), .SUM({\alu/N307 , \alu/N338 , 
        \alu/N337 , \alu/N336 , \alu/N335 , \alu/N334 , \alu/N333 , \alu/N332 , 
        \alu/N331 , \alu/N330 , \alu/N329 , \alu/N328 , \alu/N327 , \alu/N326 , 
        \alu/N293 , \alu/N292 , \alu/N291 , \alu/N290 , \alu/N289 , \alu/N288 , 
        \alu/N287 , \alu/N286 , \alu/N285 , \alu/N284 , \alu/N283 , \alu/N282 , 
        \alu/N281 }) );
  CVP14_DW_rash_2 \alu/srl_136_C23  ( .A({\alu/N88 , op2[9:0], \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* }), .DATA_TC(\*Logic0* ), .SH({n215, n216, n217, 
        n218, n219}), .SH_TC(\*Logic0* ), .B({\alu/N226 , \alu/N225 , 
        \alu/N224 , \alu/N223 , \alu/N222 , \alu/N221 , \alu/N220 , \alu/N219 , 
        \alu/N218 , \alu/N217 , \alu/N216 , \alu/N215 , \alu/N214 , \alu/N213 , 
        \alu/N212 , \alu/N211 , \alu/N210 , \alu/N209 , \alu/N208 , \alu/N207 , 
        \alu/N206 , \alu/N205 , \alu/N204 , \alu/N203 , \alu/N202 , \alu/N201 }) );
  CVP14_DW_rash_3 \alu/srl_130_C23  ( .A({\alu/N87 , op1[9:0], \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* }), .DATA_TC(\*Logic0* ), .SH({n215, n216, n217, 
        n218, n219}), .SH_TC(\*Logic0* ), .B({\alu/N117 , \alu/N116 , 
        \alu/N115 , \alu/N114 , \alu/N113 , \alu/N112 , \alu/N111 , \alu/N110 , 
        \alu/N109 , \alu/N108 , \alu/N107 , \alu/N106 , \alu/N105 , \alu/N104 , 
        \alu/N103 , \alu/N102 , \alu/N101 , \alu/N100 , \alu/N99 , \alu/N98 , 
        \alu/N97 , \alu/N96 , \alu/N95 , \alu/N94 , \alu/N93 , \alu/N92 }) );
  CVP14_DW01_addsub_7 r149 ( .A({\*Logic0* , \U3/U29/Z_4 , \U3/U29/Z_3 , 
        \U3/U29/Z_2 , \U3/U29/Z_1 , \U3/U29/Z_0 }), .B({\*Logic0* , 
        \U3/U30/Z_4 , \U3/U30/Z_3 , \U3/U30/Z_2 , \U3/U30/Z_1 , \U3/U30/Z_0 }), 
        .CI(\U3/U31/Z_0 ), .ADD_SUB(\U3/U32/Z_0 ), .SUM({n214, n215, n216, 
        n217, n218, n219}) );
  CVP14_DW01_decode_2 C1681 ( .A(cycles), .B({SYNOPSYS_UNCONNECTED__64, 
        SYNOPSYS_UNCONNECTED__65, SYNOPSYS_UNCONNECTED__66, 
        SYNOPSYS_UNCONNECTED__67, SYNOPSYS_UNCONNECTED__68, 
        SYNOPSYS_UNCONNECTED__69, SYNOPSYS_UNCONNECTED__70, 
        SYNOPSYS_UNCONNECTED__71, SYNOPSYS_UNCONNECTED__72, 
        SYNOPSYS_UNCONNECTED__73, SYNOPSYS_UNCONNECTED__74, 
        SYNOPSYS_UNCONNECTED__75, SYNOPSYS_UNCONNECTED__76, 
        SYNOPSYS_UNCONNECTED__77, SYNOPSYS_UNCONNECTED__78, 
        SYNOPSYS_UNCONNECTED__79, SYNOPSYS_UNCONNECTED__80, N1786, N1785, 
        N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, 
        N1774, N1773, N1772}) );
  CVP14_DW02_mult_0 r160 ( .A({\alu/*Logic1* , op1[9:0]}), .B({\alu/*Logic1* , 
        op2[9:0]}), .TC(\*Logic0* ), .PRODUCT({\alu/N850 , \alu/N849 , 
        \alu/N848 , \alu/N847 , \alu/N846 , \alu/N845 , \alu/N844 , \alu/N843 , 
        \alu/N842 , \alu/N841 , \alu/N840 , \alu/N839 , 
        SYNOPSYS_UNCONNECTED__81, SYNOPSYS_UNCONNECTED__82, 
        SYNOPSYS_UNCONNECTED__83, SYNOPSYS_UNCONNECTED__84, 
        SYNOPSYS_UNCONNECTED__85, SYNOPSYS_UNCONNECTED__86, 
        SYNOPSYS_UNCONNECTED__87, SYNOPSYS_UNCONNECTED__88, 
        SYNOPSYS_UNCONNECTED__89, SYNOPSYS_UNCONNECTED__90}) );
  DFQD1BWP \state_reg[3]  ( .D(N140), .CP(Clk1), .Q(state[3]) );
  DFQD1BWP \state_reg[1]  ( .D(N138), .CP(Clk1), .Q(state[1]) );
  DFQD1BWP \state_reg[0]  ( .D(N137), .CP(Clk1), .Q(state[0]) );
  DFQD1BWP \state_reg[2]  ( .D(N139), .CP(Clk1), .Q(state[2]) );
  LHD1BWP \nextInstrAddr_reg[0]  ( .E(N4047), .D(N4048), .QN(n3424) );
  LHD1BWP \nextInstrAddr_reg[4]  ( .E(N4047), .D(N4052), .QN(n3420) );
  LHD1BWP \nextInstrAddr_reg[3]  ( .E(N4047), .D(N4051), .QN(n3421) );
  LHD1BWP \nextInstrAddr_reg[2]  ( .E(N4047), .D(N4050), .QN(n3422) );
  LHD1BWP \nextInstrAddr_reg[1]  ( .E(N4047), .D(N4049), .QN(n3423) );
  LHD1BWP \nextInstrAddr_reg[5]  ( .E(N4047), .D(N4053), .QN(n3402) );
  LHD1BWP \nextInstrAddr_reg[6]  ( .E(N4047), .D(N4054), .QN(n3401) );
  LHD1BWP \nextInstrAddr_reg[7]  ( .E(N4047), .D(N4055), .QN(n3400) );
  LHD1BWP \nextInstrAddr_reg[8]  ( .E(N4047), .D(N4056), .QN(n3399) );
  LHD1BWP \nextInstrAddr_reg[9]  ( .E(N4047), .D(N4057), .QN(n3398) );
  LHD1BWP \nextInstrAddr_reg[10]  ( .E(N4047), .D(N4058), .QN(n3397) );
  LHD1BWP \nextInstrAddr_reg[11]  ( .E(N4047), .D(N4059), .QN(n3396) );
  LHD1BWP \nextInstrAddr_reg[12]  ( .E(N4047), .D(N4060), .QN(n3395) );
  LHD1BWP \nextInstrAddr_reg[13]  ( .E(N4047), .D(N4061), .QN(n3394) );
  LHD1BWP \nextInstrAddr_reg[14]  ( .E(N4047), .D(N4062), .QN(n3393) );
  LHD1BWP \nextInstrAddr_reg[15]  ( .E(N4047), .D(N4063), .QN(n3392) );
  LHD1BWP \vectorToLoad_reg[0]  ( .E(N4105), .D(N4106), .QN(n3418) );
  LHD1BWP \vectorToLoad_reg[1]  ( .E(N4105), .D(N4107), .QN(n3417) );
  LHD1BWP \vectorToLoad_reg[2]  ( .E(N4105), .D(N4108), .QN(n3416) );
  LHD1BWP \vectorToLoad_reg[3]  ( .E(N4105), .D(N4109), .QN(n3415) );
  LHD1BWP \vectorToLoad_reg[4]  ( .E(N4105), .D(N4110), .QN(n3414) );
  LHD1BWP \vectorToLoad_reg[5]  ( .E(N4105), .D(N4111), .QN(n3413) );
  LHD1BWP \vectorToLoad_reg[6]  ( .E(N4105), .D(N4112), .QN(n3412) );
  LHD1BWP \vectorToLoad_reg[7]  ( .E(N4105), .D(N4113), .QN(n3411) );
  LHD1BWP \vectorToLoad_reg[8]  ( .E(N4105), .D(N4114), .QN(n3410) );
  LHD1BWP \vectorToLoad_reg[9]  ( .E(N4105), .D(N4115), .QN(n3409) );
  LHD1BWP \vectorToLoad_reg[10]  ( .E(N4105), .D(N4116), .QN(n3408) );
  LHD1BWP \vectorToLoad_reg[11]  ( .E(N4105), .D(N4117), .QN(n3407) );
  LHD1BWP \vectorToLoad_reg[12]  ( .E(N4105), .D(N4118), .QN(n3406) );
  LHD1BWP \vectorToLoad_reg[13]  ( .E(N4105), .D(N4119), .QN(n3405) );
  LHD1BWP \vectorToLoad_reg[14]  ( .E(N4105), .D(N4120), .QN(n3404) );
  LHD1BWP \vectorToLoad_reg[15]  ( .E(N4105), .D(N4121), .QN(n3403) );
  LHD1BWP \vectorToLoad_reg[16]  ( .E(n5394), .D(N4123), .QN(n3419) );
  LHQD1BWP \memAddr_reg[1]  ( .E(N4028), .D(N4030), .Q(Addr[1]) );
  LHQD1BWP \memAddr_reg[2]  ( .E(N4028), .D(N4031), .Q(Addr[2]) );
  LHQD1BWP \memAddr_reg[3]  ( .E(N4028), .D(N4032), .Q(Addr[3]) );
  LHQD1BWP \memAddr_reg[4]  ( .E(N4028), .D(N4033), .Q(Addr[4]) );
  LHQD1BWP \memAddr_reg[5]  ( .E(N4028), .D(N4034), .Q(Addr[5]) );
  LHQD1BWP \memAddr_reg[6]  ( .E(N4028), .D(N4035), .Q(Addr[6]) );
  LHQD1BWP \memAddr_reg[7]  ( .E(N4028), .D(N4036), .Q(Addr[7]) );
  LHQD1BWP \memAddr_reg[8]  ( .E(N4028), .D(N4037), .Q(Addr[8]) );
  LHQD1BWP \memAddr_reg[9]  ( .E(N4028), .D(N4038), .Q(Addr[9]) );
  LHQD1BWP \memAddr_reg[10]  ( .E(N4028), .D(N4039), .Q(Addr[10]) );
  LHQD1BWP \memAddr_reg[11]  ( .E(N4028), .D(N4040), .Q(Addr[11]) );
  LHQD1BWP \memAddr_reg[12]  ( .E(N4028), .D(N4041), .Q(Addr[12]) );
  LHQD1BWP \memAddr_reg[13]  ( .E(N4028), .D(N4042), .Q(Addr[13]) );
  LHQD1BWP \memAddr_reg[14]  ( .E(N4028), .D(N4043), .Q(Addr[14]) );
  LHQD1BWP \memAddr_reg[15]  ( .E(N4028), .D(N4044), .Q(Addr[15]) );
  LHQD1BWP \memAddr_reg[0]  ( .E(N4028), .D(N4029), .Q(Addr[0]) );
  LHD1BWP \vectorToLoad_reg[17]  ( .E(n5381), .D(N4124), .Q(n7435) );
  LHD1BWP \vectorToLoad_reg[18]  ( .E(n5381), .D(N4125), .Q(n7434) );
  LHD1BWP \vectorToLoad_reg[19]  ( .E(n5381), .D(N4126), .Q(n7433) );
  LHD1BWP \vectorToLoad_reg[20]  ( .E(n5381), .D(N4127), .Q(n7432) );
  LHD1BWP \vectorToLoad_reg[21]  ( .E(n5381), .D(N4128), .Q(n7431) );
  LHD1BWP \vectorToLoad_reg[22]  ( .E(n5381), .D(N4129), .Q(n7430) );
  LHD1BWP \vectorToLoad_reg[23]  ( .E(n5381), .D(N4130), .Q(n7429) );
  LHD1BWP \vectorToLoad_reg[24]  ( .E(n5381), .D(N4131), .Q(n7428) );
  LHD1BWP \vectorToLoad_reg[25]  ( .E(n5381), .D(N4132), .Q(n7427) );
  LHD1BWP \vectorToLoad_reg[26]  ( .E(n5381), .D(N4133), .Q(n7426) );
  LHD1BWP \vectorToLoad_reg[27]  ( .E(n5381), .D(N4134), .Q(n7425) );
  LHD1BWP \vectorToLoad_reg[28]  ( .E(n5380), .D(N4135), .Q(n7424) );
  LHD1BWP \vectorToLoad_reg[29]  ( .E(n5380), .D(N4136), .Q(n7423) );
  LHD1BWP \vectorToLoad_reg[30]  ( .E(n5380), .D(N4137), .Q(n7422) );
  LHD1BWP \vectorToLoad_reg[31]  ( .E(n5380), .D(N4138), .Q(n7421) );
  LHD1BWP \vectorToLoad_reg[32]  ( .E(n5380), .D(N4139), .Q(n7420) );
  LHD1BWP \vectorToLoad_reg[33]  ( .E(n5380), .D(N4140), .Q(n7419) );
  LHD1BWP \vectorToLoad_reg[34]  ( .E(n5380), .D(N4141), .Q(n7418) );
  LHD1BWP \vectorToLoad_reg[35]  ( .E(n5380), .D(N4142), .Q(n7417) );
  LHD1BWP \vectorToLoad_reg[36]  ( .E(n5380), .D(N4143), .Q(n7416) );
  LHD1BWP \vectorToLoad_reg[37]  ( .E(n5380), .D(N4144), .Q(n7415) );
  LHD1BWP \vectorToLoad_reg[38]  ( .E(n5380), .D(N4145), .Q(n7414) );
  LHD1BWP \vectorToLoad_reg[39]  ( .E(n5380), .D(N4146), .Q(n7413) );
  LHD1BWP \vectorToLoad_reg[40]  ( .E(n5379), .D(N4147), .Q(n7412) );
  LHD1BWP \vectorToLoad_reg[41]  ( .E(n5379), .D(N4148), .Q(n7411) );
  LHD1BWP \vectorToLoad_reg[42]  ( .E(n5379), .D(N4149), .Q(n7410) );
  LHD1BWP \vectorToLoad_reg[43]  ( .E(n5379), .D(N4150), .Q(n7409) );
  LHD1BWP \vectorToLoad_reg[44]  ( .E(n5379), .D(N4151), .Q(n7408) );
  LHD1BWP \vectorToLoad_reg[45]  ( .E(n5379), .D(N4152), .Q(n7407) );
  LHD1BWP \vectorToLoad_reg[46]  ( .E(n5379), .D(N4153), .Q(n7406) );
  LHD1BWP \vectorToLoad_reg[47]  ( .E(n5379), .D(N4154), .Q(n7405) );
  LHD1BWP \vectorToLoad_reg[48]  ( .E(n5379), .D(N4155), .Q(n7404) );
  LHD1BWP \vectorToLoad_reg[49]  ( .E(n5379), .D(N4156), .Q(n7403) );
  LHD1BWP \vectorToLoad_reg[50]  ( .E(n5379), .D(N4157), .Q(n7402) );
  LHD1BWP \vectorToLoad_reg[51]  ( .E(n5379), .D(N4158), .Q(n7401) );
  LHD1BWP \vectorToLoad_reg[52]  ( .E(n5378), .D(N4159), .Q(n7400) );
  LHD1BWP \vectorToLoad_reg[53]  ( .E(n5378), .D(N4160), .Q(n7399) );
  LHD1BWP \vectorToLoad_reg[54]  ( .E(n5378), .D(N4161), .Q(n7398) );
  LHD1BWP \vectorToLoad_reg[55]  ( .E(n5378), .D(N4162), .Q(n7397) );
  LHD1BWP \vectorToLoad_reg[56]  ( .E(n5378), .D(N4163), .Q(n7396) );
  LHD1BWP \vectorToLoad_reg[57]  ( .E(n5378), .D(N4164), .Q(n7395) );
  LHD1BWP \vectorToLoad_reg[58]  ( .E(n5378), .D(N4165), .Q(n7394) );
  LHD1BWP \vectorToLoad_reg[59]  ( .E(n5378), .D(N4166), .Q(n7393) );
  LHD1BWP \vectorToLoad_reg[60]  ( .E(n5378), .D(N4167), .Q(n7392) );
  LHD1BWP \vectorToLoad_reg[61]  ( .E(n5378), .D(N4168), .Q(n7391) );
  LHD1BWP \vectorToLoad_reg[62]  ( .E(n5378), .D(N4169), .Q(n7390) );
  LHD1BWP \vectorToLoad_reg[63]  ( .E(n5378), .D(N4170), .Q(n7389) );
  LHD1BWP \vectorToLoad_reg[64]  ( .E(n5377), .D(N4171), .Q(n7388) );
  LHD1BWP \vectorToLoad_reg[65]  ( .E(n5377), .D(N4172), .Q(n7387) );
  LHD1BWP \vectorToLoad_reg[66]  ( .E(n5377), .D(N4173), .Q(n7386) );
  LHD1BWP \vectorToLoad_reg[67]  ( .E(n5377), .D(N4174), .Q(n7385) );
  LHD1BWP \vectorToLoad_reg[68]  ( .E(n5377), .D(N4175), .Q(n7384) );
  LHD1BWP \vectorToLoad_reg[69]  ( .E(n5377), .D(N4176), .Q(n7383) );
  LHD1BWP \vectorToLoad_reg[70]  ( .E(n5377), .D(N4177), .Q(n7382) );
  LHD1BWP \vectorToLoad_reg[71]  ( .E(n5377), .D(N4178), .Q(n7381) );
  LHD1BWP \vectorToLoad_reg[72]  ( .E(n5377), .D(N4179), .Q(n7380) );
  LHD1BWP \vectorToLoad_reg[73]  ( .E(n5377), .D(N4180), .Q(n7379) );
  LHD1BWP \vectorToLoad_reg[74]  ( .E(n5377), .D(N4181), .Q(n7378) );
  LHD1BWP \vectorToLoad_reg[75]  ( .E(n5377), .D(N4182), .Q(n7377) );
  LHD1BWP \vectorToLoad_reg[76]  ( .E(n5376), .D(N4183), .Q(n7376) );
  LHD1BWP \vectorToLoad_reg[77]  ( .E(n5376), .D(N4184), .Q(n7375) );
  LHD1BWP \vectorToLoad_reg[78]  ( .E(n5376), .D(N4185), .Q(n7374) );
  LHD1BWP \vectorToLoad_reg[79]  ( .E(n5376), .D(N4186), .Q(n7373) );
  LHD1BWP \vectorToLoad_reg[80]  ( .E(n5376), .D(N4187), .Q(n7372) );
  LHD1BWP \vectorToLoad_reg[81]  ( .E(n5376), .D(N4188), .Q(n7371) );
  LHD1BWP \vectorToLoad_reg[82]  ( .E(n5376), .D(N4189), .Q(n7370) );
  LHD1BWP \vectorToLoad_reg[83]  ( .E(n5376), .D(N4190), .Q(n7369) );
  LHD1BWP \vectorToLoad_reg[84]  ( .E(n5376), .D(N4191), .Q(n7368) );
  LHD1BWP \vectorToLoad_reg[85]  ( .E(n5376), .D(N4192), .Q(n7367) );
  LHD1BWP \vectorToLoad_reg[86]  ( .E(n5376), .D(N4193), .Q(n7366) );
  LHD1BWP \vectorToLoad_reg[87]  ( .E(n5376), .D(N4194), .Q(n7365) );
  LHD1BWP \vectorToLoad_reg[88]  ( .E(n5375), .D(N4195), .Q(n7364) );
  LHD1BWP \vectorToLoad_reg[89]  ( .E(n5375), .D(N4196), .Q(n7363) );
  LHD1BWP \vectorToLoad_reg[90]  ( .E(n5375), .D(N4197), .Q(n7362) );
  LHD1BWP \vectorToLoad_reg[91]  ( .E(n5375), .D(N4198), .Q(n7361) );
  LHD1BWP \vectorToLoad_reg[92]  ( .E(n5375), .D(N4199), .Q(n7360) );
  LHD1BWP \vectorToLoad_reg[93]  ( .E(n5375), .D(N4200), .Q(n7359) );
  LHD1BWP \vectorToLoad_reg[94]  ( .E(n5375), .D(N4201), .Q(n7358) );
  LHD1BWP \vectorToLoad_reg[95]  ( .E(n5375), .D(N4202), .Q(n7357) );
  LHD1BWP \vectorToLoad_reg[96]  ( .E(n5375), .D(N4203), .Q(n7356) );
  LHD1BWP \vectorToLoad_reg[97]  ( .E(n5375), .D(N4204), .Q(n7355) );
  LHD1BWP \vectorToLoad_reg[98]  ( .E(n5375), .D(N4205), .Q(n7354) );
  LHD1BWP \vectorToLoad_reg[99]  ( .E(n5375), .D(N4206), .Q(n7353) );
  LHD1BWP \vectorToLoad_reg[100]  ( .E(n5384), .D(N4207), .Q(n7352) );
  LHD1BWP \vectorToLoad_reg[101]  ( .E(n5384), .D(N4208), .Q(n7351) );
  LHD1BWP \vectorToLoad_reg[102]  ( .E(n5384), .D(N4209), .Q(n7350) );
  LHD1BWP \vectorToLoad_reg[103]  ( .E(n5383), .D(N4210), .Q(n7349) );
  LHD1BWP \vectorToLoad_reg[104]  ( .E(n5383), .D(N4211), .Q(n7348) );
  LHD1BWP \vectorToLoad_reg[105]  ( .E(n5383), .D(N4212), .Q(n7347) );
  LHD1BWP \vectorToLoad_reg[106]  ( .E(n5383), .D(N4213), .Q(n7346) );
  LHD1BWP \vectorToLoad_reg[107]  ( .E(n5383), .D(N4214), .Q(n7345) );
  LHD1BWP \vectorToLoad_reg[108]  ( .E(n5383), .D(N4215), .Q(n7344) );
  LHD1BWP \vectorToLoad_reg[109]  ( .E(n5383), .D(N4216), .Q(n7343) );
  LHD1BWP \vectorToLoad_reg[110]  ( .E(n5383), .D(N4217), .Q(n7342) );
  LHD1BWP \vectorToLoad_reg[111]  ( .E(n5383), .D(N4218), .Q(n7341) );
  LHD1BWP \vectorToLoad_reg[112]  ( .E(n5383), .D(N4219), .Q(n7340) );
  LHD1BWP \vectorToLoad_reg[113]  ( .E(n5383), .D(N4220), .Q(n7339) );
  LHD1BWP \vectorToLoad_reg[114]  ( .E(n5383), .D(N4221), .Q(n7338) );
  LHD1BWP \vectorToLoad_reg[115]  ( .E(n5382), .D(N4223), .Q(n7337) );
  LHD1BWP \vectorToLoad_reg[116]  ( .E(n5382), .D(N4224), .Q(n7336) );
  LHD1BWP \vectorToLoad_reg[117]  ( .E(n5382), .D(N4225), .Q(n7335) );
  LHD1BWP \vectorToLoad_reg[118]  ( .E(n5382), .D(N4226), .Q(n7334) );
  LHD1BWP \vectorToLoad_reg[119]  ( .E(n5382), .D(N4227), .Q(n7333) );
  LHD1BWP \vectorToLoad_reg[120]  ( .E(n5382), .D(N4228), .Q(n7332) );
  LHD1BWP \vectorToLoad_reg[121]  ( .E(n5382), .D(N4229), .Q(n7331) );
  LHD1BWP \vectorToLoad_reg[122]  ( .E(n5382), .D(N4230), .Q(n7330) );
  LHD1BWP \vectorToLoad_reg[123]  ( .E(n5382), .D(N4231), .Q(n7329) );
  LHD1BWP \vectorToLoad_reg[124]  ( .E(n5382), .D(N4232), .Q(n7328) );
  LHD1BWP \vectorToLoad_reg[125]  ( .E(n5382), .D(N4233), .Q(n7327) );
  LHD1BWP \vectorToLoad_reg[126]  ( .E(n5382), .D(N4234), .Q(n7326) );
  LHD1BWP \vectorToLoad_reg[127]  ( .E(n5381), .D(N4235), .Q(n7325) );
  LHD1BWP \vectorToLoad_reg[128]  ( .E(n5384), .D(N4236), .Q(n7324) );
  LHD1BWP \vectorToLoad_reg[129]  ( .E(n5384), .D(N4237), .Q(n7323) );
  LHD1BWP \vectorToLoad_reg[130]  ( .E(n5384), .D(N4238), .Q(n7322) );
  LHD1BWP \vectorToLoad_reg[131]  ( .E(n5384), .D(N4239), .Q(n7321) );
  LHD1BWP \vectorToLoad_reg[132]  ( .E(n5384), .D(N4240), .Q(n7320) );
  LHD1BWP \vectorToLoad_reg[133]  ( .E(n5384), .D(N4241), .Q(n7319) );
  LHD1BWP \vectorToLoad_reg[134]  ( .E(n5384), .D(N4242), .Q(n7318) );
  LHD1BWP \vectorToLoad_reg[135]  ( .E(n5384), .D(N4243), .Q(n7317) );
  LHD1BWP \vectorToLoad_reg[136]  ( .E(n5384), .D(N4244), .Q(n7316) );
  LHD1BWP \vectorToLoad_reg[137]  ( .E(n5385), .D(N4245), .Q(n7315) );
  LHD1BWP \vectorToLoad_reg[138]  ( .E(n5385), .D(N4246), .Q(n7314) );
  LHD1BWP \vectorToLoad_reg[139]  ( .E(n5385), .D(N4247), .Q(n7313) );
  LHD1BWP \vectorToLoad_reg[140]  ( .E(n5385), .D(N4248), .Q(n7312) );
  LHD1BWP \vectorToLoad_reg[141]  ( .E(n5385), .D(N4249), .Q(n7311) );
  LHD1BWP \vectorToLoad_reg[142]  ( .E(n5385), .D(N4250), .Q(n7310) );
  LHD1BWP \vectorToLoad_reg[143]  ( .E(n5385), .D(N4251), .Q(n7309) );
  LHD1BWP \vectorToLoad_reg[144]  ( .E(n5385), .D(N4252), .Q(n7308) );
  LHD1BWP \vectorToLoad_reg[145]  ( .E(n5385), .D(N4253), .Q(n7307) );
  LHD1BWP \vectorToLoad_reg[146]  ( .E(n5385), .D(N4254), .Q(n7306) );
  LHD1BWP \vectorToLoad_reg[147]  ( .E(n5385), .D(N4255), .Q(n7305) );
  LHD1BWP \vectorToLoad_reg[148]  ( .E(n5385), .D(N4256), .Q(n7304) );
  LHD1BWP \vectorToLoad_reg[149]  ( .E(n5386), .D(N4257), .Q(n7303) );
  LHD1BWP \vectorToLoad_reg[150]  ( .E(n5386), .D(N4258), .Q(n7302) );
  LHD1BWP \vectorToLoad_reg[151]  ( .E(n5386), .D(N4259), .Q(n7301) );
  LHD1BWP \vectorToLoad_reg[152]  ( .E(n5386), .D(N4260), .Q(n7300) );
  LHD1BWP \vectorToLoad_reg[153]  ( .E(n5386), .D(N4261), .Q(n7299) );
  LHD1BWP \vectorToLoad_reg[154]  ( .E(n5386), .D(N4262), .Q(n7298) );
  LHD1BWP \vectorToLoad_reg[155]  ( .E(n5386), .D(N4263), .Q(n7297) );
  LHD1BWP \vectorToLoad_reg[156]  ( .E(n5386), .D(N4264), .Q(n7296) );
  LHD1BWP \vectorToLoad_reg[157]  ( .E(n5386), .D(N4265), .Q(n7295) );
  LHD1BWP \vectorToLoad_reg[158]  ( .E(n5386), .D(N4266), .Q(n7294) );
  LHD1BWP \vectorToLoad_reg[159]  ( .E(n5386), .D(N4267), .Q(n7293) );
  LHD1BWP \vectorToLoad_reg[160]  ( .E(n5386), .D(N4268), .Q(n7292) );
  LHD1BWP \vectorToLoad_reg[161]  ( .E(n5387), .D(N4269), .Q(n7291) );
  LHD1BWP \vectorToLoad_reg[162]  ( .E(n5387), .D(N4270), .Q(n7290) );
  LHD1BWP \vectorToLoad_reg[163]  ( .E(n5387), .D(N4271), .Q(n7289) );
  LHD1BWP \vectorToLoad_reg[164]  ( .E(n5387), .D(N4272), .Q(n7288) );
  LHD1BWP \vectorToLoad_reg[165]  ( .E(n5387), .D(N4273), .Q(n7287) );
  LHD1BWP \vectorToLoad_reg[166]  ( .E(n5387), .D(N4274), .Q(n7286) );
  LHD1BWP \vectorToLoad_reg[167]  ( .E(n5387), .D(N4275), .Q(n7285) );
  LHD1BWP \vectorToLoad_reg[168]  ( .E(n5387), .D(N4276), .Q(n7284) );
  LHD1BWP \vectorToLoad_reg[169]  ( .E(n5387), .D(N4277), .Q(n7283) );
  LHD1BWP \vectorToLoad_reg[170]  ( .E(n5387), .D(N4278), .Q(n7282) );
  LHD1BWP \vectorToLoad_reg[171]  ( .E(n5387), .D(N4279), .Q(n7281) );
  LHD1BWP \vectorToLoad_reg[172]  ( .E(n5387), .D(N4280), .Q(n7280) );
  LHD1BWP \vectorToLoad_reg[173]  ( .E(n5388), .D(N4281), .Q(n7279) );
  LHD1BWP \vectorToLoad_reg[174]  ( .E(n5388), .D(N4282), .Q(n7278) );
  LHD1BWP \vectorToLoad_reg[175]  ( .E(n5388), .D(N4283), .Q(n7277) );
  LHD1BWP \vectorToLoad_reg[176]  ( .E(n5388), .D(N4284), .Q(n7276) );
  LHD1BWP \vectorToLoad_reg[177]  ( .E(n5388), .D(N4285), .Q(n7275) );
  LHD1BWP \vectorToLoad_reg[178]  ( .E(n5388), .D(N4286), .Q(n7274) );
  LHD1BWP \vectorToLoad_reg[179]  ( .E(n5388), .D(N4287), .Q(n7273) );
  LHD1BWP \vectorToLoad_reg[180]  ( .E(n5388), .D(N4288), .Q(n7272) );
  LHD1BWP \vectorToLoad_reg[181]  ( .E(n5388), .D(N4289), .Q(n7271) );
  LHD1BWP \vectorToLoad_reg[182]  ( .E(n5388), .D(N4290), .Q(n7270) );
  LHD1BWP \vectorToLoad_reg[183]  ( .E(n5388), .D(N4291), .Q(n7269) );
  LHD1BWP \vectorToLoad_reg[184]  ( .E(n5388), .D(N4292), .Q(n7268) );
  LHD1BWP \vectorToLoad_reg[185]  ( .E(n5389), .D(N4293), .Q(n7267) );
  LHD1BWP \vectorToLoad_reg[186]  ( .E(n5389), .D(N4294), .Q(n7266) );
  LHD1BWP \vectorToLoad_reg[187]  ( .E(n5389), .D(N4295), .Q(n7265) );
  LHD1BWP \vectorToLoad_reg[188]  ( .E(n5389), .D(N4296), .Q(n7264) );
  LHD1BWP \vectorToLoad_reg[189]  ( .E(n5389), .D(N4297), .Q(n7263) );
  LHD1BWP \vectorToLoad_reg[190]  ( .E(n5389), .D(N4298), .Q(n7262) );
  LHD1BWP \vectorToLoad_reg[191]  ( .E(n5389), .D(N4299), .Q(n7261) );
  LHD1BWP \vectorToLoad_reg[192]  ( .E(n5389), .D(N4300), .Q(n7260) );
  LHD1BWP \vectorToLoad_reg[193]  ( .E(n5389), .D(N4301), .Q(n7259) );
  LHD1BWP \vectorToLoad_reg[194]  ( .E(n5389), .D(N4302), .Q(n7258) );
  LHD1BWP \vectorToLoad_reg[195]  ( .E(n5389), .D(N4303), .Q(n7257) );
  LHD1BWP \vectorToLoad_reg[196]  ( .E(n5389), .D(N4304), .Q(n7256) );
  LHD1BWP \vectorToLoad_reg[197]  ( .E(n5390), .D(N4305), .Q(n7255) );
  LHD1BWP \vectorToLoad_reg[198]  ( .E(n5390), .D(N4306), .Q(n7254) );
  LHD1BWP \vectorToLoad_reg[199]  ( .E(n5390), .D(N4307), .Q(n7253) );
  LHD1BWP \vectorToLoad_reg[200]  ( .E(n5390), .D(N4308), .Q(n7252) );
  LHD1BWP \vectorToLoad_reg[201]  ( .E(n5390), .D(N4309), .Q(n7251) );
  LHD1BWP \vectorToLoad_reg[202]  ( .E(n5390), .D(N4310), .Q(n7250) );
  LHD1BWP \vectorToLoad_reg[203]  ( .E(n5390), .D(N4311), .Q(n7249) );
  LHD1BWP \vectorToLoad_reg[204]  ( .E(n5390), .D(N4312), .Q(n7248) );
  LHD1BWP \vectorToLoad_reg[205]  ( .E(n5390), .D(N4313), .Q(n7247) );
  LHD1BWP \vectorToLoad_reg[206]  ( .E(n5390), .D(N4314), .Q(n7246) );
  LHD1BWP \vectorToLoad_reg[207]  ( .E(n5390), .D(N4315), .Q(n7245) );
  LHD1BWP \vectorToLoad_reg[208]  ( .E(n5390), .D(N4316), .Q(n7244) );
  LHD1BWP \vectorToLoad_reg[209]  ( .E(n5391), .D(N4317), .Q(n7243) );
  LHD1BWP \vectorToLoad_reg[210]  ( .E(n5391), .D(N4318), .Q(n7242) );
  LHD1BWP \vectorToLoad_reg[211]  ( .E(n5391), .D(N4319), .Q(n7241) );
  LHD1BWP \vectorToLoad_reg[212]  ( .E(n5391), .D(N4320), .Q(n7240) );
  LHD1BWP \vectorToLoad_reg[213]  ( .E(n5391), .D(N4321), .Q(n7239) );
  LHD1BWP \vectorToLoad_reg[214]  ( .E(n5391), .D(N4323), .Q(n7238) );
  LHD1BWP \vectorToLoad_reg[215]  ( .E(n5391), .D(N4324), .Q(n7237) );
  LHD1BWP \vectorToLoad_reg[216]  ( .E(n5391), .D(N4325), .Q(n7236) );
  LHD1BWP \vectorToLoad_reg[217]  ( .E(n5391), .D(N4326), .Q(n7235) );
  LHD1BWP \vectorToLoad_reg[218]  ( .E(n5391), .D(N4327), .Q(n7234) );
  LHD1BWP \vectorToLoad_reg[219]  ( .E(n5391), .D(N4328), .Q(n7233) );
  LHD1BWP \vectorToLoad_reg[220]  ( .E(n5391), .D(N4329), .Q(n7232) );
  LHD1BWP \vectorToLoad_reg[221]  ( .E(n5392), .D(N4330), .Q(n7231) );
  LHD1BWP \vectorToLoad_reg[222]  ( .E(n5392), .D(N4331), .Q(n7230) );
  LHD1BWP \vectorToLoad_reg[223]  ( .E(n5392), .D(N4332), .Q(n7229) );
  LHD1BWP \vectorToLoad_reg[224]  ( .E(n5392), .D(N4333), .Q(n7228) );
  LHD1BWP \vectorToLoad_reg[225]  ( .E(n5392), .D(N4334), .Q(n7227) );
  LHD1BWP \vectorToLoad_reg[226]  ( .E(n5392), .D(N4335), .Q(n7226) );
  LHD1BWP \vectorToLoad_reg[227]  ( .E(n5392), .D(N4336), .Q(n7225) );
  LHD1BWP \vectorToLoad_reg[228]  ( .E(n5392), .D(N4337), .Q(n7224) );
  LHD1BWP \vectorToLoad_reg[229]  ( .E(n5392), .D(N4338), .Q(n7223) );
  LHD1BWP \vectorToLoad_reg[230]  ( .E(n5392), .D(N4339), .Q(n7222) );
  LHD1BWP \vectorToLoad_reg[231]  ( .E(n5392), .D(N4340), .Q(n7221) );
  LHD1BWP \vectorToLoad_reg[232]  ( .E(n5392), .D(N4341), .Q(n7220) );
  LHD1BWP \vectorToLoad_reg[233]  ( .E(n5393), .D(N4342), .Q(n7219) );
  LHD1BWP \vectorToLoad_reg[234]  ( .E(n5393), .D(N4343), .Q(n7218) );
  LHD1BWP \vectorToLoad_reg[235]  ( .E(n5393), .D(N4344), .Q(n7217) );
  LHD1BWP \vectorToLoad_reg[236]  ( .E(n5393), .D(N4345), .Q(n7216) );
  LHD1BWP \vectorToLoad_reg[237]  ( .E(n5393), .D(N4346), .Q(n7215) );
  LHD1BWP \vectorToLoad_reg[238]  ( .E(n5393), .D(N4347), .Q(n7214) );
  LHD1BWP \vectorToLoad_reg[239]  ( .E(n5393), .D(N4348), .Q(n7213) );
  LHD1BWP \vectorToLoad_reg[240]  ( .E(n5393), .D(N4349), .Q(n7212) );
  LHD1BWP \vectorToLoad_reg[241]  ( .E(n5393), .D(N4350), .Q(n7211) );
  LHD1BWP \vectorToLoad_reg[242]  ( .E(n5393), .D(N4351), .Q(n7210) );
  LHD1BWP \vectorToLoad_reg[243]  ( .E(n5393), .D(N4352), .Q(n7209) );
  LHD1BWP \vectorToLoad_reg[244]  ( .E(n5393), .D(N4353), .Q(n7208) );
  LHD1BWP \vectorToLoad_reg[245]  ( .E(n5394), .D(N4354), .Q(n7207) );
  LHD1BWP \vectorToLoad_reg[246]  ( .E(n5394), .D(N4355), .Q(n7206) );
  LHD1BWP \vectorToLoad_reg[247]  ( .E(n5394), .D(N4356), .Q(n7205) );
  LHD1BWP \vectorToLoad_reg[248]  ( .E(n5394), .D(N4357), .Q(n7204) );
  LHD1BWP \vectorToLoad_reg[249]  ( .E(n5394), .D(N4358), .Q(n7203) );
  LHD1BWP \vectorToLoad_reg[250]  ( .E(n5394), .D(N4359), .Q(n7202) );
  LHD1BWP \vectorToLoad_reg[251]  ( .E(n5394), .D(N4360), .Q(n7201) );
  LHD1BWP \vectorToLoad_reg[252]  ( .E(n5394), .D(N4361), .Q(n7200) );
  LHD1BWP \vectorToLoad_reg[253]  ( .E(n5394), .D(N4362), .Q(n7199) );
  LHD1BWP \vectorToLoad_reg[254]  ( .E(n5394), .D(N4363), .Q(n7198) );
  LHD1BWP \vectorToLoad_reg[255]  ( .E(n5394), .D(N4364), .Q(n7197) );
  LNQD1BWP \instrIn_reg[3]  ( .D(DataIn[3]), .EN(n3262), .Q(instrIn[3]) );
  LNQD1BWP \instrIn_reg[4]  ( .D(DataIn[4]), .EN(n3262), .Q(instrIn[4]) );
  LNQD1BWP \instrIn_reg[0]  ( .D(DataIn[0]), .EN(n3262), .Q(instrIn[0]) );
  LNQD1BWP \scalarWrData_reg[10]  ( .D(N3763), .EN(n1461), .Q(scalarWrData[10]) );
  LNQD1BWP \scalarWrData_reg[14]  ( .D(N3767), .EN(n1461), .Q(scalarWrData[14]) );
  LNQD1BWP \scalarWrData_reg[13]  ( .D(N3766), .EN(n1461), .Q(scalarWrData[13]) );
  LNQD1BWP \scalarWrData_reg[12]  ( .D(N3765), .EN(n1461), .Q(scalarWrData[12]) );
  LNQD1BWP \scalarWrData_reg[11]  ( .D(N3764), .EN(n1461), .Q(scalarWrData[11]) );
  LNQD1BWP \scalarWrData_reg[15]  ( .D(N3768), .EN(n1461), .Q(scalarWrData[15]) );
  LNQD1BWP \scalarWrData_reg[9]  ( .D(N3762), .EN(n1461), .Q(scalarWrData[9])
         );
  LNQD1BWP \scalarWrData_reg[8]  ( .D(N3761), .EN(n1461), .Q(scalarWrData[8])
         );
  LNQD1BWP \scalarWrData_reg[7]  ( .D(N3760), .EN(n1461), .Q(scalarWrData[7])
         );
  LNQD1BWP \scalarWrData_reg[6]  ( .D(N3759), .EN(n1461), .Q(scalarWrData[6])
         );
  LNQD1BWP \scalarWrData_reg[5]  ( .D(N3758), .EN(n1461), .Q(scalarWrData[5])
         );
  LNQD1BWP \scalarWrData_reg[4]  ( .D(N3757), .EN(n1461), .Q(scalarWrData[4])
         );
  LNQD1BWP \scalarWrData_reg[3]  ( .D(N3756), .EN(n1461), .Q(scalarWrData[3])
         );
  LNQD1BWP \scalarWrData_reg[2]  ( .D(N3755), .EN(n1461), .Q(scalarWrData[2])
         );
  LNQD1BWP \scalarWrData_reg[1]  ( .D(N3754), .EN(n1461), .Q(scalarWrData[1])
         );
  LNQD1BWP \scalarWrData_reg[0]  ( .D(N3753), .EN(n1461), .Q(scalarWrData[0])
         );
  LNQD1BWP \instrIn_reg[1]  ( .D(DataIn[1]), .EN(n3262), .Q(instrIn[1]) );
  LNQD1BWP \instrIn_reg[2]  ( .D(DataIn[2]), .EN(n3262), .Q(instrIn[2]) );
  LHQD1BWP \wrAddr_reg[2]  ( .E(N4366), .D(addrDst[2]), .Q(\srf/N17 ) );
  LHQD1BWP \op2_reg[15]  ( .E(N4102), .D(N4101), .Q(op2[15]) );
  LNQD1BWP \instrIn_reg[11]  ( .D(DataIn[11]), .EN(n3262), .Q(instrIn[11]) );
  LNQD1BWP \instrIn_reg[5]  ( .D(DataIn[5]), .EN(n3262), .Q(instrIn[5]) );
  LNQD1BWP \instrIn_reg[6]  ( .D(DataIn[6]), .EN(n3262), .Q(instrIn[6]) );
  LNQD1BWP \instrIn_reg[7]  ( .D(DataIn[7]), .EN(n3262), .Q(instrIn[7]) );
  LNQD1BWP \instrIn_reg[8]  ( .D(DataIn[8]), .EN(n3262), .Q(instrIn[8]) );
  LNQD1BWP \instrIn_reg[9]  ( .D(DataIn[9]), .EN(n3262), .Q(instrIn[9]) );
  LNQD1BWP \instrIn_reg[10]  ( .D(DataIn[10]), .EN(n3262), .Q(instrIn[10]) );
  LHQD1BWP \op2_reg[14]  ( .E(N4102), .D(N4100), .Q(op2[14]) );
  LNQD1BWP \scalarToLoad_reg[11]  ( .D(N1758), .EN(n2522), .Q(scalarToLoad[11]) );
  LNQD1BWP \scalarToLoad_reg[15]  ( .D(N1762), .EN(n2522), .Q(scalarToLoad[15]) );
  LHQD1BWP \vrf/regTable_reg[5][15]  ( .E(n5192), .D(\vrf/N33 ), .Q(
        \vrf/regTable[5][15] ) );
  LHQD1BWP \vrf/regTable_reg[5][16]  ( .E(n5192), .D(\vrf/N34 ), .Q(
        \vrf/regTable[5][16] ) );
  LHQD1BWP \vrf/regTable_reg[5][254]  ( .E(n5192), .D(\vrf/N274 ), .Q(
        \vrf/regTable[5][254] ) );
  LHQD1BWP \vrf/regTable_reg[5][255]  ( .E(n5192), .D(\vrf/N275 ), .Q(
        \vrf/regTable[5][255] ) );
  LHQD1BWP \vrf/regTable_reg[1][15]  ( .E(n5328), .D(\vrf/N33 ), .Q(
        \vrf/regTable[1][15] ) );
  LHQD1BWP \vrf/regTable_reg[1][16]  ( .E(n5328), .D(\vrf/N34 ), .Q(
        \vrf/regTable[1][16] ) );
  LHQD1BWP \vrf/regTable_reg[1][254]  ( .E(n5328), .D(\vrf/N274 ), .Q(
        \vrf/regTable[1][254] ) );
  LHQD1BWP \vrf/regTable_reg[1][255]  ( .E(n5328), .D(\vrf/N275 ), .Q(
        \vrf/regTable[1][255] ) );
  LHQD1BWP \vrf/regTable_reg[5][0]  ( .E(n5181), .D(\vrf/N18 ), .Q(
        \vrf/regTable[5][0] ) );
  LHQD1BWP \vrf/regTable_reg[5][1]  ( .E(n5178), .D(\vrf/N19 ), .Q(
        \vrf/regTable[5][1] ) );
  LHQD1BWP \vrf/regTable_reg[5][2]  ( .E(n5177), .D(\vrf/N20 ), .Q(
        \vrf/regTable[5][2] ) );
  LHQD1BWP \vrf/regTable_reg[5][3]  ( .E(n5176), .D(\vrf/N21 ), .Q(
        \vrf/regTable[5][3] ) );
  LHQD1BWP \vrf/regTable_reg[5][4]  ( .E(n5175), .D(\vrf/N22 ), .Q(
        \vrf/regTable[5][4] ) );
  LHQD1BWP \vrf/regTable_reg[5][5]  ( .E(n5174), .D(\vrf/N23 ), .Q(
        \vrf/regTable[5][5] ) );
  LHQD1BWP \vrf/regTable_reg[5][6]  ( .E(n5173), .D(\vrf/N24 ), .Q(
        \vrf/regTable[5][6] ) );
  LHQD1BWP \vrf/regTable_reg[5][7]  ( .E(n5172), .D(\vrf/N25 ), .Q(
        \vrf/regTable[5][7] ) );
  LHQD1BWP \vrf/regTable_reg[5][8]  ( .E(n5171), .D(\vrf/N26 ), .Q(
        \vrf/regTable[5][8] ) );
  LHQD1BWP \vrf/regTable_reg[5][9]  ( .E(n5171), .D(\vrf/N27 ), .Q(
        \vrf/regTable[5][9] ) );
  LHQD1BWP \vrf/regTable_reg[5][10]  ( .E(n5180), .D(\vrf/N28 ), .Q(
        \vrf/regTable[5][10] ) );
  LHQD1BWP \vrf/regTable_reg[5][11]  ( .E(n5179), .D(\vrf/N29 ), .Q(
        \vrf/regTable[5][11] ) );
  LHQD1BWP \vrf/regTable_reg[5][12]  ( .E(n5178), .D(\vrf/N30 ), .Q(
        \vrf/regTable[5][12] ) );
  LHQD1BWP \vrf/regTable_reg[5][13]  ( .E(n5178), .D(\vrf/N31 ), .Q(
        \vrf/regTable[5][13] ) );
  LHQD1BWP \vrf/regTable_reg[5][14]  ( .E(n5178), .D(\vrf/N32 ), .Q(
        \vrf/regTable[5][14] ) );
  LHQD1BWP \vrf/regTable_reg[5][17]  ( .E(n5178), .D(\vrf/N35 ), .Q(
        \vrf/regTable[5][17] ) );
  LHQD1BWP \vrf/regTable_reg[5][18]  ( .E(n5178), .D(\vrf/N36 ), .Q(
        \vrf/regTable[5][18] ) );
  LHQD1BWP \vrf/regTable_reg[5][19]  ( .E(n5178), .D(\vrf/N37 ), .Q(
        \vrf/regTable[5][19] ) );
  LHQD1BWP \vrf/regTable_reg[5][20]  ( .E(n5178), .D(\vrf/N38 ), .Q(
        \vrf/regTable[5][20] ) );
  LHQD1BWP \vrf/regTable_reg[5][21]  ( .E(n5178), .D(\vrf/N39 ), .Q(
        \vrf/regTable[5][21] ) );
  LHQD1BWP \vrf/regTable_reg[5][22]  ( .E(n5178), .D(\vrf/N40 ), .Q(
        \vrf/regTable[5][22] ) );
  LHQD1BWP \vrf/regTable_reg[5][23]  ( .E(n5178), .D(\vrf/N41 ), .Q(
        \vrf/regTable[5][23] ) );
  LHQD1BWP \vrf/regTable_reg[5][24]  ( .E(n5177), .D(\vrf/N42 ), .Q(
        \vrf/regTable[5][24] ) );
  LHQD1BWP \vrf/regTable_reg[5][25]  ( .E(n5177), .D(\vrf/N43 ), .Q(
        \vrf/regTable[5][25] ) );
  LHQD1BWP \vrf/regTable_reg[5][26]  ( .E(n5177), .D(\vrf/N44 ), .Q(
        \vrf/regTable[5][26] ) );
  LHQD1BWP \vrf/regTable_reg[5][27]  ( .E(n5177), .D(\vrf/N45 ), .Q(
        \vrf/regTable[5][27] ) );
  LHQD1BWP \vrf/regTable_reg[5][28]  ( .E(n5177), .D(\vrf/N46 ), .Q(
        \vrf/regTable[5][28] ) );
  LHQD1BWP \vrf/regTable_reg[5][29]  ( .E(n5177), .D(\vrf/N47 ), .Q(
        \vrf/regTable[5][29] ) );
  LHQD1BWP \vrf/regTable_reg[5][30]  ( .E(n5177), .D(\vrf/N48 ), .Q(
        \vrf/regTable[5][30] ) );
  LHQD1BWP \vrf/regTable_reg[5][31]  ( .E(n5177), .D(\vrf/N49 ), .Q(
        \vrf/regTable[5][31] ) );
  LHQD1BWP \vrf/regTable_reg[5][32]  ( .E(n5177), .D(\vrf/N50 ), .Q(
        \vrf/regTable[5][32] ) );
  LHQD1BWP \vrf/regTable_reg[5][33]  ( .E(n5177), .D(\vrf/N51 ), .Q(
        \vrf/regTable[5][33] ) );
  LHQD1BWP \vrf/regTable_reg[5][34]  ( .E(n5177), .D(\vrf/N52 ), .Q(
        \vrf/regTable[5][34] ) );
  LHQD1BWP \vrf/regTable_reg[5][35]  ( .E(n5176), .D(\vrf/N53 ), .Q(
        \vrf/regTable[5][35] ) );
  LHQD1BWP \vrf/regTable_reg[5][36]  ( .E(n5176), .D(\vrf/N54 ), .Q(
        \vrf/regTable[5][36] ) );
  LHQD1BWP \vrf/regTable_reg[5][37]  ( .E(n5176), .D(\vrf/N55 ), .Q(
        \vrf/regTable[5][37] ) );
  LHQD1BWP \vrf/regTable_reg[5][38]  ( .E(n5176), .D(\vrf/N56 ), .Q(
        \vrf/regTable[5][38] ) );
  LHQD1BWP \vrf/regTable_reg[5][39]  ( .E(n5176), .D(\vrf/N57 ), .Q(
        \vrf/regTable[5][39] ) );
  LHQD1BWP \vrf/regTable_reg[5][40]  ( .E(n5176), .D(\vrf/N58 ), .Q(
        \vrf/regTable[5][40] ) );
  LHQD1BWP \vrf/regTable_reg[5][41]  ( .E(n5176), .D(\vrf/N59 ), .Q(
        \vrf/regTable[5][41] ) );
  LHQD1BWP \vrf/regTable_reg[5][42]  ( .E(n5176), .D(\vrf/N60 ), .Q(
        \vrf/regTable[5][42] ) );
  LHQD1BWP \vrf/regTable_reg[5][43]  ( .E(n5176), .D(\vrf/N61 ), .Q(
        \vrf/regTable[5][43] ) );
  LHQD1BWP \vrf/regTable_reg[5][44]  ( .E(n5176), .D(\vrf/N62 ), .Q(
        \vrf/regTable[5][44] ) );
  LHQD1BWP \vrf/regTable_reg[5][45]  ( .E(n5176), .D(\vrf/N63 ), .Q(
        \vrf/regTable[5][45] ) );
  LHQD1BWP \vrf/regTable_reg[5][46]  ( .E(n5175), .D(\vrf/N64 ), .Q(
        \vrf/regTable[5][46] ) );
  LHQD1BWP \vrf/regTable_reg[5][47]  ( .E(n5175), .D(\vrf/N65 ), .Q(
        \vrf/regTable[5][47] ) );
  LHQD1BWP \vrf/regTable_reg[5][48]  ( .E(n5175), .D(\vrf/N66 ), .Q(
        \vrf/regTable[5][48] ) );
  LHQD1BWP \vrf/regTable_reg[5][49]  ( .E(n5175), .D(\vrf/N67 ), .Q(
        \vrf/regTable[5][49] ) );
  LHQD1BWP \vrf/regTable_reg[5][50]  ( .E(n5175), .D(\vrf/N68 ), .Q(
        \vrf/regTable[5][50] ) );
  LHQD1BWP \vrf/regTable_reg[5][51]  ( .E(n5175), .D(\vrf/N69 ), .Q(
        \vrf/regTable[5][51] ) );
  LHQD1BWP \vrf/regTable_reg[5][52]  ( .E(n5175), .D(\vrf/N70 ), .Q(
        \vrf/regTable[5][52] ) );
  LHQD1BWP \vrf/regTable_reg[5][53]  ( .E(n5175), .D(\vrf/N71 ), .Q(
        \vrf/regTable[5][53] ) );
  LHQD1BWP \vrf/regTable_reg[5][54]  ( .E(n5175), .D(\vrf/N72 ), .Q(
        \vrf/regTable[5][54] ) );
  LHQD1BWP \vrf/regTable_reg[5][55]  ( .E(n5175), .D(\vrf/N73 ), .Q(
        \vrf/regTable[5][55] ) );
  LHQD1BWP \vrf/regTable_reg[5][56]  ( .E(n5175), .D(\vrf/N74 ), .Q(
        \vrf/regTable[5][56] ) );
  LHQD1BWP \vrf/regTable_reg[5][57]  ( .E(n5174), .D(\vrf/N75 ), .Q(
        \vrf/regTable[5][57] ) );
  LHQD1BWP \vrf/regTable_reg[5][58]  ( .E(n5174), .D(\vrf/N76 ), .Q(
        \vrf/regTable[5][58] ) );
  LHQD1BWP \vrf/regTable_reg[5][59]  ( .E(n5174), .D(\vrf/N77 ), .Q(
        \vrf/regTable[5][59] ) );
  LHQD1BWP \vrf/regTable_reg[5][60]  ( .E(n5174), .D(\vrf/N78 ), .Q(
        \vrf/regTable[5][60] ) );
  LHQD1BWP \vrf/regTable_reg[5][61]  ( .E(n5174), .D(\vrf/N79 ), .Q(
        \vrf/regTable[5][61] ) );
  LHQD1BWP \vrf/regTable_reg[5][62]  ( .E(n5174), .D(\vrf/N80 ), .Q(
        \vrf/regTable[5][62] ) );
  LHQD1BWP \vrf/regTable_reg[5][63]  ( .E(n5174), .D(\vrf/N81 ), .Q(
        \vrf/regTable[5][63] ) );
  LHQD1BWP \vrf/regTable_reg[5][64]  ( .E(n5174), .D(\vrf/N82 ), .Q(
        \vrf/regTable[5][64] ) );
  LHQD1BWP \vrf/regTable_reg[5][65]  ( .E(n5174), .D(\vrf/N83 ), .Q(
        \vrf/regTable[5][65] ) );
  LHQD1BWP \vrf/regTable_reg[5][66]  ( .E(n5174), .D(\vrf/N84 ), .Q(
        \vrf/regTable[5][66] ) );
  LHQD1BWP \vrf/regTable_reg[5][67]  ( .E(n5174), .D(\vrf/N85 ), .Q(
        \vrf/regTable[5][67] ) );
  LHQD1BWP \vrf/regTable_reg[5][68]  ( .E(n5173), .D(\vrf/N86 ), .Q(
        \vrf/regTable[5][68] ) );
  LHQD1BWP \vrf/regTable_reg[5][69]  ( .E(n5173), .D(\vrf/N87 ), .Q(
        \vrf/regTable[5][69] ) );
  LHQD1BWP \vrf/regTable_reg[5][70]  ( .E(n5173), .D(\vrf/N88 ), .Q(
        \vrf/regTable[5][70] ) );
  LHQD1BWP \vrf/regTable_reg[5][71]  ( .E(n5173), .D(\vrf/N89 ), .Q(
        \vrf/regTable[5][71] ) );
  LHQD1BWP \vrf/regTable_reg[5][72]  ( .E(n5173), .D(\vrf/N90 ), .Q(
        \vrf/regTable[5][72] ) );
  LHQD1BWP \vrf/regTable_reg[5][73]  ( .E(n5173), .D(\vrf/N91 ), .Q(
        \vrf/regTable[5][73] ) );
  LHQD1BWP \vrf/regTable_reg[5][74]  ( .E(n5173), .D(\vrf/N92 ), .Q(
        \vrf/regTable[5][74] ) );
  LHQD1BWP \vrf/regTable_reg[5][75]  ( .E(n5173), .D(\vrf/N93 ), .Q(
        \vrf/regTable[5][75] ) );
  LHQD1BWP \vrf/regTable_reg[5][76]  ( .E(n5173), .D(\vrf/N94 ), .Q(
        \vrf/regTable[5][76] ) );
  LHQD1BWP \vrf/regTable_reg[5][77]  ( .E(n5173), .D(\vrf/N95 ), .Q(
        \vrf/regTable[5][77] ) );
  LHQD1BWP \vrf/regTable_reg[5][78]  ( .E(n5173), .D(\vrf/N96 ), .Q(
        \vrf/regTable[5][78] ) );
  LHQD1BWP \vrf/regTable_reg[5][79]  ( .E(n5172), .D(\vrf/N97 ), .Q(
        \vrf/regTable[5][79] ) );
  LHQD1BWP \vrf/regTable_reg[5][80]  ( .E(n5172), .D(\vrf/N98 ), .Q(
        \vrf/regTable[5][80] ) );
  LHQD1BWP \vrf/regTable_reg[5][81]  ( .E(n5172), .D(\vrf/N99 ), .Q(
        \vrf/regTable[5][81] ) );
  LHQD1BWP \vrf/regTable_reg[5][82]  ( .E(n5172), .D(\vrf/N100 ), .Q(
        \vrf/regTable[5][82] ) );
  LHQD1BWP \vrf/regTable_reg[5][83]  ( .E(n5172), .D(\vrf/N101 ), .Q(
        \vrf/regTable[5][83] ) );
  LHQD1BWP \vrf/regTable_reg[5][84]  ( .E(n5172), .D(\vrf/N102 ), .Q(
        \vrf/regTable[5][84] ) );
  LHQD1BWP \vrf/regTable_reg[5][85]  ( .E(n5172), .D(\vrf/N103 ), .Q(
        \vrf/regTable[5][85] ) );
  LHQD1BWP \vrf/regTable_reg[5][86]  ( .E(n5172), .D(\vrf/N104 ), .Q(
        \vrf/regTable[5][86] ) );
  LHQD1BWP \vrf/regTable_reg[5][87]  ( .E(n5172), .D(\vrf/N105 ), .Q(
        \vrf/regTable[5][87] ) );
  LHQD1BWP \vrf/regTable_reg[5][88]  ( .E(n5172), .D(\vrf/N106 ), .Q(
        \vrf/regTable[5][88] ) );
  LHQD1BWP \vrf/regTable_reg[5][89]  ( .E(n5172), .D(\vrf/N107 ), .Q(
        \vrf/regTable[5][89] ) );
  LHQD1BWP \vrf/regTable_reg[5][90]  ( .E(n5171), .D(\vrf/N108 ), .Q(
        \vrf/regTable[5][90] ) );
  LHQD1BWP \vrf/regTable_reg[5][91]  ( .E(n5171), .D(\vrf/N109 ), .Q(
        \vrf/regTable[5][91] ) );
  LHQD1BWP \vrf/regTable_reg[5][92]  ( .E(n5171), .D(\vrf/N110 ), .Q(
        \vrf/regTable[5][92] ) );
  LHQD1BWP \vrf/regTable_reg[5][93]  ( .E(n5171), .D(\vrf/N111 ), .Q(
        \vrf/regTable[5][93] ) );
  LHQD1BWP \vrf/regTable_reg[5][94]  ( .E(n5171), .D(\vrf/N112 ), .Q(
        \vrf/regTable[5][94] ) );
  LHQD1BWP \vrf/regTable_reg[5][95]  ( .E(n5171), .D(\vrf/N113 ), .Q(
        \vrf/regTable[5][95] ) );
  LHQD1BWP \vrf/regTable_reg[5][96]  ( .E(n5171), .D(\vrf/N114 ), .Q(
        \vrf/regTable[5][96] ) );
  LHQD1BWP \vrf/regTable_reg[5][97]  ( .E(n5171), .D(\vrf/N115 ), .Q(
        \vrf/regTable[5][97] ) );
  LHQD1BWP \vrf/regTable_reg[5][98]  ( .E(n5171), .D(\vrf/N116 ), .Q(
        \vrf/regTable[5][98] ) );
  LHQD1BWP \vrf/regTable_reg[5][99]  ( .E(n5171), .D(\vrf/N118 ), .Q(
        \vrf/regTable[5][99] ) );
  LHQD1BWP \vrf/regTable_reg[5][100]  ( .E(n5181), .D(\vrf/N119 ), .Q(
        \vrf/regTable[5][100] ) );
  LHQD1BWP \vrf/regTable_reg[5][101]  ( .E(n5181), .D(\vrf/N120 ), .Q(
        \vrf/regTable[5][101] ) );
  LHQD1BWP \vrf/regTable_reg[5][102]  ( .E(n5181), .D(\vrf/N121 ), .Q(
        \vrf/regTable[5][102] ) );
  LHQD1BWP \vrf/regTable_reg[5][103]  ( .E(n5181), .D(\vrf/N122 ), .Q(
        \vrf/regTable[5][103] ) );
  LHQD1BWP \vrf/regTable_reg[5][104]  ( .E(n5181), .D(\vrf/N123 ), .Q(
        \vrf/regTable[5][104] ) );
  LHQD1BWP \vrf/regTable_reg[5][105]  ( .E(n5180), .D(\vrf/N124 ), .Q(
        \vrf/regTable[5][105] ) );
  LHQD1BWP \vrf/regTable_reg[5][106]  ( .E(n5180), .D(\vrf/N125 ), .Q(
        \vrf/regTable[5][106] ) );
  LHQD1BWP \vrf/regTable_reg[5][107]  ( .E(n5180), .D(\vrf/N126 ), .Q(
        \vrf/regTable[5][107] ) );
  LHQD1BWP \vrf/regTable_reg[5][108]  ( .E(n5180), .D(\vrf/N127 ), .Q(
        \vrf/regTable[5][108] ) );
  LHQD1BWP \vrf/regTable_reg[5][109]  ( .E(n5180), .D(\vrf/N128 ), .Q(
        \vrf/regTable[5][109] ) );
  LHQD1BWP \vrf/regTable_reg[5][110]  ( .E(n5180), .D(\vrf/N129 ), .Q(
        \vrf/regTable[5][110] ) );
  LHQD1BWP \vrf/regTable_reg[5][111]  ( .E(n5180), .D(\vrf/N130 ), .Q(
        \vrf/regTable[5][111] ) );
  LHQD1BWP \vrf/regTable_reg[5][112]  ( .E(n5180), .D(\vrf/N131 ), .Q(
        \vrf/regTable[5][112] ) );
  LHQD1BWP \vrf/regTable_reg[5][113]  ( .E(n5180), .D(\vrf/N132 ), .Q(
        \vrf/regTable[5][113] ) );
  LHQD1BWP \vrf/regTable_reg[5][114]  ( .E(n5180), .D(\vrf/N133 ), .Q(
        \vrf/regTable[5][114] ) );
  LHQD1BWP \vrf/regTable_reg[5][115]  ( .E(n5180), .D(\vrf/N134 ), .Q(
        \vrf/regTable[5][115] ) );
  LHQD1BWP \vrf/regTable_reg[5][116]  ( .E(n5179), .D(\vrf/N135 ), .Q(
        \vrf/regTable[5][116] ) );
  LHQD1BWP \vrf/regTable_reg[5][117]  ( .E(n5179), .D(\vrf/N136 ), .Q(
        \vrf/regTable[5][117] ) );
  LHQD1BWP \vrf/regTable_reg[5][118]  ( .E(n5179), .D(\vrf/N137 ), .Q(
        \vrf/regTable[5][118] ) );
  LHQD1BWP \vrf/regTable_reg[5][119]  ( .E(n5179), .D(\vrf/N138 ), .Q(
        \vrf/regTable[5][119] ) );
  LHQD1BWP \vrf/regTable_reg[5][120]  ( .E(n5179), .D(\vrf/N139 ), .Q(
        \vrf/regTable[5][120] ) );
  LHQD1BWP \vrf/regTable_reg[5][121]  ( .E(n5179), .D(\vrf/N140 ), .Q(
        \vrf/regTable[5][121] ) );
  LHQD1BWP \vrf/regTable_reg[5][122]  ( .E(n5179), .D(\vrf/N141 ), .Q(
        \vrf/regTable[5][122] ) );
  LHQD1BWP \vrf/regTable_reg[5][123]  ( .E(n5179), .D(\vrf/N142 ), .Q(
        \vrf/regTable[5][123] ) );
  LHQD1BWP \vrf/regTable_reg[5][124]  ( .E(n5179), .D(\vrf/N143 ), .Q(
        \vrf/regTable[5][124] ) );
  LHQD1BWP \vrf/regTable_reg[5][125]  ( .E(n5179), .D(\vrf/N144 ), .Q(
        \vrf/regTable[5][125] ) );
  LHQD1BWP \vrf/regTable_reg[5][126]  ( .E(n5179), .D(\vrf/N145 ), .Q(
        \vrf/regTable[5][126] ) );
  LHQD1BWP \vrf/regTable_reg[5][127]  ( .E(n5178), .D(\vrf/N146 ), .Q(
        \vrf/regTable[5][127] ) );
  LHQD1BWP \vrf/regTable_reg[5][128]  ( .E(n5181), .D(\vrf/N147 ), .Q(
        \vrf/regTable[5][128] ) );
  LHQD1BWP \vrf/regTable_reg[5][129]  ( .E(n5181), .D(\vrf/N148 ), .Q(
        \vrf/regTable[5][129] ) );
  LHQD1BWP \vrf/regTable_reg[5][130]  ( .E(n5181), .D(\vrf/N149 ), .Q(
        \vrf/regTable[5][130] ) );
  LHQD1BWP \vrf/regTable_reg[5][131]  ( .E(n5181), .D(\vrf/N150 ), .Q(
        \vrf/regTable[5][131] ) );
  LHQD1BWP \vrf/regTable_reg[5][132]  ( .E(n5181), .D(\vrf/N151 ), .Q(
        \vrf/regTable[5][132] ) );
  LHQD1BWP \vrf/regTable_reg[5][133]  ( .E(n5181), .D(\vrf/N152 ), .Q(
        \vrf/regTable[5][133] ) );
  LHQD1BWP \vrf/regTable_reg[5][134]  ( .E(n5182), .D(\vrf/N153 ), .Q(
        \vrf/regTable[5][134] ) );
  LHQD1BWP \vrf/regTable_reg[5][135]  ( .E(n5182), .D(\vrf/N154 ), .Q(
        \vrf/regTable[5][135] ) );
  LHQD1BWP \vrf/regTable_reg[5][136]  ( .E(n5182), .D(\vrf/N155 ), .Q(
        \vrf/regTable[5][136] ) );
  LHQD1BWP \vrf/regTable_reg[5][137]  ( .E(n5182), .D(\vrf/N156 ), .Q(
        \vrf/regTable[5][137] ) );
  LHQD1BWP \vrf/regTable_reg[5][138]  ( .E(n5182), .D(\vrf/N157 ), .Q(
        \vrf/regTable[5][138] ) );
  LHQD1BWP \vrf/regTable_reg[5][139]  ( .E(n5182), .D(\vrf/N158 ), .Q(
        \vrf/regTable[5][139] ) );
  LHQD1BWP \vrf/regTable_reg[5][140]  ( .E(n5182), .D(\vrf/N159 ), .Q(
        \vrf/regTable[5][140] ) );
  LHQD1BWP \vrf/regTable_reg[5][141]  ( .E(n5182), .D(\vrf/N160 ), .Q(
        \vrf/regTable[5][141] ) );
  LHQD1BWP \vrf/regTable_reg[5][142]  ( .E(n5182), .D(\vrf/N161 ), .Q(
        \vrf/regTable[5][142] ) );
  LHQD1BWP \vrf/regTable_reg[5][143]  ( .E(n5182), .D(\vrf/N162 ), .Q(
        \vrf/regTable[5][143] ) );
  LHQD1BWP \vrf/regTable_reg[5][144]  ( .E(n5182), .D(\vrf/N163 ), .Q(
        \vrf/regTable[5][144] ) );
  LHQD1BWP \vrf/regTable_reg[5][145]  ( .E(n5182), .D(\vrf/N164 ), .Q(
        \vrf/regTable[5][145] ) );
  LHQD1BWP \vrf/regTable_reg[5][146]  ( .E(n5183), .D(\vrf/N165 ), .Q(
        \vrf/regTable[5][146] ) );
  LHQD1BWP \vrf/regTable_reg[5][147]  ( .E(n5183), .D(\vrf/N166 ), .Q(
        \vrf/regTable[5][147] ) );
  LHQD1BWP \vrf/regTable_reg[5][148]  ( .E(n5183), .D(\vrf/N167 ), .Q(
        \vrf/regTable[5][148] ) );
  LHQD1BWP \vrf/regTable_reg[5][149]  ( .E(n5183), .D(\vrf/N168 ), .Q(
        \vrf/regTable[5][149] ) );
  LHQD1BWP \vrf/regTable_reg[5][150]  ( .E(n5183), .D(\vrf/N169 ), .Q(
        \vrf/regTable[5][150] ) );
  LHQD1BWP \vrf/regTable_reg[5][151]  ( .E(n5183), .D(\vrf/N170 ), .Q(
        \vrf/regTable[5][151] ) );
  LHQD1BWP \vrf/regTable_reg[5][152]  ( .E(n5183), .D(\vrf/N171 ), .Q(
        \vrf/regTable[5][152] ) );
  LHQD1BWP \vrf/regTable_reg[5][153]  ( .E(n5183), .D(\vrf/N172 ), .Q(
        \vrf/regTable[5][153] ) );
  LHQD1BWP \vrf/regTable_reg[5][154]  ( .E(n5183), .D(\vrf/N173 ), .Q(
        \vrf/regTable[5][154] ) );
  LHQD1BWP \vrf/regTable_reg[5][155]  ( .E(n5183), .D(\vrf/N174 ), .Q(
        \vrf/regTable[5][155] ) );
  LHQD1BWP \vrf/regTable_reg[5][156]  ( .E(n5183), .D(\vrf/N175 ), .Q(
        \vrf/regTable[5][156] ) );
  LHQD1BWP \vrf/regTable_reg[5][157]  ( .E(n5183), .D(\vrf/N176 ), .Q(
        \vrf/regTable[5][157] ) );
  LHQD1BWP \vrf/regTable_reg[5][158]  ( .E(n5184), .D(\vrf/N177 ), .Q(
        \vrf/regTable[5][158] ) );
  LHQD1BWP \vrf/regTable_reg[5][159]  ( .E(n5184), .D(\vrf/N178 ), .Q(
        \vrf/regTable[5][159] ) );
  LHQD1BWP \vrf/regTable_reg[5][160]  ( .E(n5184), .D(\vrf/N179 ), .Q(
        \vrf/regTable[5][160] ) );
  LHQD1BWP \vrf/regTable_reg[5][161]  ( .E(n5184), .D(\vrf/N180 ), .Q(
        \vrf/regTable[5][161] ) );
  LHQD1BWP \vrf/regTable_reg[5][162]  ( .E(n5184), .D(\vrf/N181 ), .Q(
        \vrf/regTable[5][162] ) );
  LHQD1BWP \vrf/regTable_reg[5][163]  ( .E(n5184), .D(\vrf/N182 ), .Q(
        \vrf/regTable[5][163] ) );
  LHQD1BWP \vrf/regTable_reg[5][164]  ( .E(n5184), .D(\vrf/N183 ), .Q(
        \vrf/regTable[5][164] ) );
  LHQD1BWP \vrf/regTable_reg[5][165]  ( .E(n5184), .D(\vrf/N184 ), .Q(
        \vrf/regTable[5][165] ) );
  LHQD1BWP \vrf/regTable_reg[5][166]  ( .E(n5184), .D(\vrf/N185 ), .Q(
        \vrf/regTable[5][166] ) );
  LHQD1BWP \vrf/regTable_reg[5][167]  ( .E(n5184), .D(\vrf/N186 ), .Q(
        \vrf/regTable[5][167] ) );
  LHQD1BWP \vrf/regTable_reg[5][168]  ( .E(n5184), .D(\vrf/N187 ), .Q(
        \vrf/regTable[5][168] ) );
  LHQD1BWP \vrf/regTable_reg[5][169]  ( .E(n5184), .D(\vrf/N188 ), .Q(
        \vrf/regTable[5][169] ) );
  LHQD1BWP \vrf/regTable_reg[5][170]  ( .E(n5185), .D(\vrf/N189 ), .Q(
        \vrf/regTable[5][170] ) );
  LHQD1BWP \vrf/regTable_reg[5][171]  ( .E(n5185), .D(\vrf/N190 ), .Q(
        \vrf/regTable[5][171] ) );
  LHQD1BWP \vrf/regTable_reg[5][172]  ( .E(n5185), .D(\vrf/N191 ), .Q(
        \vrf/regTable[5][172] ) );
  LHQD1BWP \vrf/regTable_reg[5][173]  ( .E(n5185), .D(\vrf/N192 ), .Q(
        \vrf/regTable[5][173] ) );
  LHQD1BWP \vrf/regTable_reg[5][174]  ( .E(n5185), .D(\vrf/N193 ), .Q(
        \vrf/regTable[5][174] ) );
  LHQD1BWP \vrf/regTable_reg[5][175]  ( .E(n5185), .D(\vrf/N194 ), .Q(
        \vrf/regTable[5][175] ) );
  LHQD1BWP \vrf/regTable_reg[5][176]  ( .E(n5185), .D(\vrf/N195 ), .Q(
        \vrf/regTable[5][176] ) );
  LHQD1BWP \vrf/regTable_reg[5][177]  ( .E(n5185), .D(\vrf/N196 ), .Q(
        \vrf/regTable[5][177] ) );
  LHQD1BWP \vrf/regTable_reg[5][178]  ( .E(n5185), .D(\vrf/N197 ), .Q(
        \vrf/regTable[5][178] ) );
  LHQD1BWP \vrf/regTable_reg[5][179]  ( .E(n5185), .D(\vrf/N198 ), .Q(
        \vrf/regTable[5][179] ) );
  LHQD1BWP \vrf/regTable_reg[5][180]  ( .E(n5185), .D(\vrf/N199 ), .Q(
        \vrf/regTable[5][180] ) );
  LHQD1BWP \vrf/regTable_reg[5][181]  ( .E(n5185), .D(\vrf/N200 ), .Q(
        \vrf/regTable[5][181] ) );
  LHQD1BWP \vrf/regTable_reg[5][182]  ( .E(n5186), .D(\vrf/N201 ), .Q(
        \vrf/regTable[5][182] ) );
  LHQD1BWP \vrf/regTable_reg[5][183]  ( .E(n5186), .D(\vrf/N202 ), .Q(
        \vrf/regTable[5][183] ) );
  LHQD1BWP \vrf/regTable_reg[5][184]  ( .E(n5186), .D(\vrf/N203 ), .Q(
        \vrf/regTable[5][184] ) );
  LHQD1BWP \vrf/regTable_reg[5][185]  ( .E(n5186), .D(\vrf/N204 ), .Q(
        \vrf/regTable[5][185] ) );
  LHQD1BWP \vrf/regTable_reg[5][186]  ( .E(n5186), .D(\vrf/N205 ), .Q(
        \vrf/regTable[5][186] ) );
  LHQD1BWP \vrf/regTable_reg[5][187]  ( .E(n5186), .D(\vrf/N206 ), .Q(
        \vrf/regTable[5][187] ) );
  LHQD1BWP \vrf/regTable_reg[5][188]  ( .E(n5186), .D(\vrf/N207 ), .Q(
        \vrf/regTable[5][188] ) );
  LHQD1BWP \vrf/regTable_reg[5][189]  ( .E(n5186), .D(\vrf/N208 ), .Q(
        \vrf/regTable[5][189] ) );
  LHQD1BWP \vrf/regTable_reg[5][190]  ( .E(n5186), .D(\vrf/N209 ), .Q(
        \vrf/regTable[5][190] ) );
  LHQD1BWP \vrf/regTable_reg[5][191]  ( .E(n5186), .D(\vrf/N210 ), .Q(
        \vrf/regTable[5][191] ) );
  LHQD1BWP \vrf/regTable_reg[5][192]  ( .E(n5186), .D(\vrf/N211 ), .Q(
        \vrf/regTable[5][192] ) );
  LHQD1BWP \vrf/regTable_reg[5][193]  ( .E(n5186), .D(\vrf/N212 ), .Q(
        \vrf/regTable[5][193] ) );
  LHQD1BWP \vrf/regTable_reg[5][194]  ( .E(n5187), .D(\vrf/N213 ), .Q(
        \vrf/regTable[5][194] ) );
  LHQD1BWP \vrf/regTable_reg[5][195]  ( .E(n5187), .D(\vrf/N214 ), .Q(
        \vrf/regTable[5][195] ) );
  LHQD1BWP \vrf/regTable_reg[5][196]  ( .E(n5187), .D(\vrf/N215 ), .Q(
        \vrf/regTable[5][196] ) );
  LHQD1BWP \vrf/regTable_reg[5][197]  ( .E(n5187), .D(\vrf/N216 ), .Q(
        \vrf/regTable[5][197] ) );
  LHQD1BWP \vrf/regTable_reg[5][198]  ( .E(n5187), .D(\vrf/N218 ), .Q(
        \vrf/regTable[5][198] ) );
  LHQD1BWP \vrf/regTable_reg[5][199]  ( .E(n5187), .D(\vrf/N219 ), .Q(
        \vrf/regTable[5][199] ) );
  LHQD1BWP \vrf/regTable_reg[5][200]  ( .E(n5187), .D(\vrf/N220 ), .Q(
        \vrf/regTable[5][200] ) );
  LHQD1BWP \vrf/regTable_reg[5][201]  ( .E(n5187), .D(\vrf/N221 ), .Q(
        \vrf/regTable[5][201] ) );
  LHQD1BWP \vrf/regTable_reg[5][202]  ( .E(n5187), .D(\vrf/N222 ), .Q(
        \vrf/regTable[5][202] ) );
  LHQD1BWP \vrf/regTable_reg[5][203]  ( .E(n5187), .D(\vrf/N223 ), .Q(
        \vrf/regTable[5][203] ) );
  LHQD1BWP \vrf/regTable_reg[5][204]  ( .E(n5187), .D(\vrf/N224 ), .Q(
        \vrf/regTable[5][204] ) );
  LHQD1BWP \vrf/regTable_reg[5][205]  ( .E(n5187), .D(\vrf/N225 ), .Q(
        \vrf/regTable[5][205] ) );
  LHQD1BWP \vrf/regTable_reg[5][206]  ( .E(n5188), .D(\vrf/N226 ), .Q(
        \vrf/regTable[5][206] ) );
  LHQD1BWP \vrf/regTable_reg[5][207]  ( .E(n5188), .D(\vrf/N227 ), .Q(
        \vrf/regTable[5][207] ) );
  LHQD1BWP \vrf/regTable_reg[5][208]  ( .E(n5188), .D(\vrf/N228 ), .Q(
        \vrf/regTable[5][208] ) );
  LHQD1BWP \vrf/regTable_reg[5][209]  ( .E(n5188), .D(\vrf/N229 ), .Q(
        \vrf/regTable[5][209] ) );
  LHQD1BWP \vrf/regTable_reg[5][210]  ( .E(n5188), .D(\vrf/N230 ), .Q(
        \vrf/regTable[5][210] ) );
  LHQD1BWP \vrf/regTable_reg[5][211]  ( .E(n5188), .D(\vrf/N231 ), .Q(
        \vrf/regTable[5][211] ) );
  LHQD1BWP \vrf/regTable_reg[5][212]  ( .E(n5188), .D(\vrf/N232 ), .Q(
        \vrf/regTable[5][212] ) );
  LHQD1BWP \vrf/regTable_reg[5][213]  ( .E(n5188), .D(\vrf/N233 ), .Q(
        \vrf/regTable[5][213] ) );
  LHQD1BWP \vrf/regTable_reg[5][214]  ( .E(n5188), .D(\vrf/N234 ), .Q(
        \vrf/regTable[5][214] ) );
  LHQD1BWP \vrf/regTable_reg[5][215]  ( .E(n5188), .D(\vrf/N235 ), .Q(
        \vrf/regTable[5][215] ) );
  LHQD1BWP \vrf/regTable_reg[5][216]  ( .E(n5188), .D(\vrf/N236 ), .Q(
        \vrf/regTable[5][216] ) );
  LHQD1BWP \vrf/regTable_reg[5][217]  ( .E(n5188), .D(\vrf/N237 ), .Q(
        \vrf/regTable[5][217] ) );
  LHQD1BWP \vrf/regTable_reg[5][218]  ( .E(n5189), .D(\vrf/N238 ), .Q(
        \vrf/regTable[5][218] ) );
  LHQD1BWP \vrf/regTable_reg[5][219]  ( .E(n5189), .D(\vrf/N239 ), .Q(
        \vrf/regTable[5][219] ) );
  LHQD1BWP \vrf/regTable_reg[5][220]  ( .E(n5189), .D(\vrf/N240 ), .Q(
        \vrf/regTable[5][220] ) );
  LHQD1BWP \vrf/regTable_reg[5][221]  ( .E(n5189), .D(\vrf/N241 ), .Q(
        \vrf/regTable[5][221] ) );
  LHQD1BWP \vrf/regTable_reg[5][222]  ( .E(n5189), .D(\vrf/N242 ), .Q(
        \vrf/regTable[5][222] ) );
  LHQD1BWP \vrf/regTable_reg[5][223]  ( .E(n5189), .D(\vrf/N243 ), .Q(
        \vrf/regTable[5][223] ) );
  LHQD1BWP \vrf/regTable_reg[5][224]  ( .E(n5189), .D(\vrf/N244 ), .Q(
        \vrf/regTable[5][224] ) );
  LHQD1BWP \vrf/regTable_reg[5][225]  ( .E(n5189), .D(\vrf/N245 ), .Q(
        \vrf/regTable[5][225] ) );
  LHQD1BWP \vrf/regTable_reg[5][226]  ( .E(n5189), .D(\vrf/N246 ), .Q(
        \vrf/regTable[5][226] ) );
  LHQD1BWP \vrf/regTable_reg[5][227]  ( .E(n5189), .D(\vrf/N247 ), .Q(
        \vrf/regTable[5][227] ) );
  LHQD1BWP \vrf/regTable_reg[5][228]  ( .E(n5189), .D(\vrf/N248 ), .Q(
        \vrf/regTable[5][228] ) );
  LHQD1BWP \vrf/regTable_reg[5][229]  ( .E(n5189), .D(\vrf/N249 ), .Q(
        \vrf/regTable[5][229] ) );
  LHQD1BWP \vrf/regTable_reg[5][230]  ( .E(n5190), .D(\vrf/N250 ), .Q(
        \vrf/regTable[5][230] ) );
  LHQD1BWP \vrf/regTable_reg[5][231]  ( .E(n5190), .D(\vrf/N251 ), .Q(
        \vrf/regTable[5][231] ) );
  LHQD1BWP \vrf/regTable_reg[5][232]  ( .E(n5190), .D(\vrf/N252 ), .Q(
        \vrf/regTable[5][232] ) );
  LHQD1BWP \vrf/regTable_reg[5][233]  ( .E(n5190), .D(\vrf/N253 ), .Q(
        \vrf/regTable[5][233] ) );
  LHQD1BWP \vrf/regTable_reg[5][234]  ( .E(n5190), .D(\vrf/N254 ), .Q(
        \vrf/regTable[5][234] ) );
  LHQD1BWP \vrf/regTable_reg[5][235]  ( .E(n5190), .D(\vrf/N255 ), .Q(
        \vrf/regTable[5][235] ) );
  LHQD1BWP \vrf/regTable_reg[5][236]  ( .E(n5190), .D(\vrf/N256 ), .Q(
        \vrf/regTable[5][236] ) );
  LHQD1BWP \vrf/regTable_reg[5][237]  ( .E(n5190), .D(\vrf/N257 ), .Q(
        \vrf/regTable[5][237] ) );
  LHQD1BWP \vrf/regTable_reg[5][238]  ( .E(n5190), .D(\vrf/N258 ), .Q(
        \vrf/regTable[5][238] ) );
  LHQD1BWP \vrf/regTable_reg[5][239]  ( .E(n5190), .D(\vrf/N259 ), .Q(
        \vrf/regTable[5][239] ) );
  LHQD1BWP \vrf/regTable_reg[5][240]  ( .E(n5190), .D(\vrf/N260 ), .Q(
        \vrf/regTable[5][240] ) );
  LHQD1BWP \vrf/regTable_reg[5][241]  ( .E(n5190), .D(\vrf/N261 ), .Q(
        \vrf/regTable[5][241] ) );
  LHQD1BWP \vrf/regTable_reg[5][242]  ( .E(n5191), .D(\vrf/N262 ), .Q(
        \vrf/regTable[5][242] ) );
  LHQD1BWP \vrf/regTable_reg[5][243]  ( .E(n5191), .D(\vrf/N263 ), .Q(
        \vrf/regTable[5][243] ) );
  LHQD1BWP \vrf/regTable_reg[5][244]  ( .E(n5191), .D(\vrf/N264 ), .Q(
        \vrf/regTable[5][244] ) );
  LHQD1BWP \vrf/regTable_reg[5][245]  ( .E(n5191), .D(\vrf/N265 ), .Q(
        \vrf/regTable[5][245] ) );
  LHQD1BWP \vrf/regTable_reg[5][246]  ( .E(n5191), .D(\vrf/N266 ), .Q(
        \vrf/regTable[5][246] ) );
  LHQD1BWP \vrf/regTable_reg[5][247]  ( .E(n5191), .D(\vrf/N267 ), .Q(
        \vrf/regTable[5][247] ) );
  LHQD1BWP \vrf/regTable_reg[5][248]  ( .E(n5191), .D(\vrf/N268 ), .Q(
        \vrf/regTable[5][248] ) );
  LHQD1BWP \vrf/regTable_reg[5][249]  ( .E(n5191), .D(\vrf/N269 ), .Q(
        \vrf/regTable[5][249] ) );
  LHQD1BWP \vrf/regTable_reg[5][250]  ( .E(n5191), .D(\vrf/N270 ), .Q(
        \vrf/regTable[5][250] ) );
  LHQD1BWP \vrf/regTable_reg[5][251]  ( .E(n5191), .D(\vrf/N271 ), .Q(
        \vrf/regTable[5][251] ) );
  LHQD1BWP \vrf/regTable_reg[5][252]  ( .E(n5191), .D(\vrf/N272 ), .Q(
        \vrf/regTable[5][252] ) );
  LHQD1BWP \vrf/regTable_reg[5][253]  ( .E(n5191), .D(\vrf/N273 ), .Q(
        \vrf/regTable[5][253] ) );
  LHQD1BWP \vrf/regTable_reg[1][0]  ( .E(n5317), .D(\vrf/N18 ), .Q(
        \vrf/regTable[1][0] ) );
  LHQD1BWP \vrf/regTable_reg[1][1]  ( .E(n5314), .D(\vrf/N19 ), .Q(
        \vrf/regTable[1][1] ) );
  LHQD1BWP \vrf/regTable_reg[1][2]  ( .E(n5313), .D(\vrf/N20 ), .Q(
        \vrf/regTable[1][2] ) );
  LHQD1BWP \vrf/regTable_reg[1][3]  ( .E(n5312), .D(\vrf/N21 ), .Q(
        \vrf/regTable[1][3] ) );
  LHQD1BWP \vrf/regTable_reg[1][4]  ( .E(n5311), .D(\vrf/N22 ), .Q(
        \vrf/regTable[1][4] ) );
  LHQD1BWP \vrf/regTable_reg[1][5]  ( .E(n5310), .D(\vrf/N23 ), .Q(
        \vrf/regTable[1][5] ) );
  LHQD1BWP \vrf/regTable_reg[1][6]  ( .E(n5309), .D(\vrf/N24 ), .Q(
        \vrf/regTable[1][6] ) );
  LHQD1BWP \vrf/regTable_reg[1][7]  ( .E(n5308), .D(\vrf/N25 ), .Q(
        \vrf/regTable[1][7] ) );
  LHQD1BWP \vrf/regTable_reg[1][8]  ( .E(n5307), .D(\vrf/N26 ), .Q(
        \vrf/regTable[1][8] ) );
  LHQD1BWP \vrf/regTable_reg[1][9]  ( .E(n5307), .D(\vrf/N27 ), .Q(
        \vrf/regTable[1][9] ) );
  LHQD1BWP \vrf/regTable_reg[1][10]  ( .E(n5316), .D(\vrf/N28 ), .Q(
        \vrf/regTable[1][10] ) );
  LHQD1BWP \vrf/regTable_reg[1][11]  ( .E(n5315), .D(\vrf/N29 ), .Q(
        \vrf/regTable[1][11] ) );
  LHQD1BWP \vrf/regTable_reg[1][12]  ( .E(n5314), .D(\vrf/N30 ), .Q(
        \vrf/regTable[1][12] ) );
  LHQD1BWP \vrf/regTable_reg[1][13]  ( .E(n5314), .D(\vrf/N31 ), .Q(
        \vrf/regTable[1][13] ) );
  LHQD1BWP \vrf/regTable_reg[1][14]  ( .E(n5314), .D(\vrf/N32 ), .Q(
        \vrf/regTable[1][14] ) );
  LHQD1BWP \vrf/regTable_reg[1][17]  ( .E(n5314), .D(\vrf/N35 ), .Q(
        \vrf/regTable[1][17] ) );
  LHQD1BWP \vrf/regTable_reg[1][18]  ( .E(n5314), .D(\vrf/N36 ), .Q(
        \vrf/regTable[1][18] ) );
  LHQD1BWP \vrf/regTable_reg[1][19]  ( .E(n5314), .D(\vrf/N37 ), .Q(
        \vrf/regTable[1][19] ) );
  LHQD1BWP \vrf/regTable_reg[1][20]  ( .E(n5314), .D(\vrf/N38 ), .Q(
        \vrf/regTable[1][20] ) );
  LHQD1BWP \vrf/regTable_reg[1][21]  ( .E(n5314), .D(\vrf/N39 ), .Q(
        \vrf/regTable[1][21] ) );
  LHQD1BWP \vrf/regTable_reg[1][22]  ( .E(n5314), .D(\vrf/N40 ), .Q(
        \vrf/regTable[1][22] ) );
  LHQD1BWP \vrf/regTable_reg[1][23]  ( .E(n5314), .D(\vrf/N41 ), .Q(
        \vrf/regTable[1][23] ) );
  LHQD1BWP \vrf/regTable_reg[1][24]  ( .E(n5313), .D(\vrf/N42 ), .Q(
        \vrf/regTable[1][24] ) );
  LHQD1BWP \vrf/regTable_reg[1][25]  ( .E(n5313), .D(\vrf/N43 ), .Q(
        \vrf/regTable[1][25] ) );
  LHQD1BWP \vrf/regTable_reg[1][26]  ( .E(n5313), .D(\vrf/N44 ), .Q(
        \vrf/regTable[1][26] ) );
  LHQD1BWP \vrf/regTable_reg[1][27]  ( .E(n5313), .D(\vrf/N45 ), .Q(
        \vrf/regTable[1][27] ) );
  LHQD1BWP \vrf/regTable_reg[1][28]  ( .E(n5313), .D(\vrf/N46 ), .Q(
        \vrf/regTable[1][28] ) );
  LHQD1BWP \vrf/regTable_reg[1][29]  ( .E(n5313), .D(\vrf/N47 ), .Q(
        \vrf/regTable[1][29] ) );
  LHQD1BWP \vrf/regTable_reg[1][30]  ( .E(n5313), .D(\vrf/N48 ), .Q(
        \vrf/regTable[1][30] ) );
  LHQD1BWP \vrf/regTable_reg[1][31]  ( .E(n5313), .D(\vrf/N49 ), .Q(
        \vrf/regTable[1][31] ) );
  LHQD1BWP \vrf/regTable_reg[1][32]  ( .E(n5313), .D(\vrf/N50 ), .Q(
        \vrf/regTable[1][32] ) );
  LHQD1BWP \vrf/regTable_reg[1][33]  ( .E(n5313), .D(\vrf/N51 ), .Q(
        \vrf/regTable[1][33] ) );
  LHQD1BWP \vrf/regTable_reg[1][34]  ( .E(n5313), .D(\vrf/N52 ), .Q(
        \vrf/regTable[1][34] ) );
  LHQD1BWP \vrf/regTable_reg[1][35]  ( .E(n5312), .D(\vrf/N53 ), .Q(
        \vrf/regTable[1][35] ) );
  LHQD1BWP \vrf/regTable_reg[1][36]  ( .E(n5312), .D(\vrf/N54 ), .Q(
        \vrf/regTable[1][36] ) );
  LHQD1BWP \vrf/regTable_reg[1][37]  ( .E(n5312), .D(\vrf/N55 ), .Q(
        \vrf/regTable[1][37] ) );
  LHQD1BWP \vrf/regTable_reg[1][38]  ( .E(n5312), .D(\vrf/N56 ), .Q(
        \vrf/regTable[1][38] ) );
  LHQD1BWP \vrf/regTable_reg[1][39]  ( .E(n5312), .D(\vrf/N57 ), .Q(
        \vrf/regTable[1][39] ) );
  LHQD1BWP \vrf/regTable_reg[1][40]  ( .E(n5312), .D(\vrf/N58 ), .Q(
        \vrf/regTable[1][40] ) );
  LHQD1BWP \vrf/regTable_reg[1][41]  ( .E(n5312), .D(\vrf/N59 ), .Q(
        \vrf/regTable[1][41] ) );
  LHQD1BWP \vrf/regTable_reg[1][42]  ( .E(n5312), .D(\vrf/N60 ), .Q(
        \vrf/regTable[1][42] ) );
  LHQD1BWP \vrf/regTable_reg[1][43]  ( .E(n5312), .D(\vrf/N61 ), .Q(
        \vrf/regTable[1][43] ) );
  LHQD1BWP \vrf/regTable_reg[1][44]  ( .E(n5312), .D(\vrf/N62 ), .Q(
        \vrf/regTable[1][44] ) );
  LHQD1BWP \vrf/regTable_reg[1][45]  ( .E(n5312), .D(\vrf/N63 ), .Q(
        \vrf/regTable[1][45] ) );
  LHQD1BWP \vrf/regTable_reg[1][46]  ( .E(n5311), .D(\vrf/N64 ), .Q(
        \vrf/regTable[1][46] ) );
  LHQD1BWP \vrf/regTable_reg[1][47]  ( .E(n5311), .D(\vrf/N65 ), .Q(
        \vrf/regTable[1][47] ) );
  LHQD1BWP \vrf/regTable_reg[1][48]  ( .E(n5311), .D(\vrf/N66 ), .Q(
        \vrf/regTable[1][48] ) );
  LHQD1BWP \vrf/regTable_reg[1][49]  ( .E(n5311), .D(\vrf/N67 ), .Q(
        \vrf/regTable[1][49] ) );
  LHQD1BWP \vrf/regTable_reg[1][50]  ( .E(n5311), .D(\vrf/N68 ), .Q(
        \vrf/regTable[1][50] ) );
  LHQD1BWP \vrf/regTable_reg[1][51]  ( .E(n5311), .D(\vrf/N69 ), .Q(
        \vrf/regTable[1][51] ) );
  LHQD1BWP \vrf/regTable_reg[1][52]  ( .E(n5311), .D(\vrf/N70 ), .Q(
        \vrf/regTable[1][52] ) );
  LHQD1BWP \vrf/regTable_reg[1][53]  ( .E(n5311), .D(\vrf/N71 ), .Q(
        \vrf/regTable[1][53] ) );
  LHQD1BWP \vrf/regTable_reg[1][54]  ( .E(n5311), .D(\vrf/N72 ), .Q(
        \vrf/regTable[1][54] ) );
  LHQD1BWP \vrf/regTable_reg[1][55]  ( .E(n5311), .D(\vrf/N73 ), .Q(
        \vrf/regTable[1][55] ) );
  LHQD1BWP \vrf/regTable_reg[1][56]  ( .E(n5311), .D(\vrf/N74 ), .Q(
        \vrf/regTable[1][56] ) );
  LHQD1BWP \vrf/regTable_reg[1][57]  ( .E(n5310), .D(\vrf/N75 ), .Q(
        \vrf/regTable[1][57] ) );
  LHQD1BWP \vrf/regTable_reg[1][58]  ( .E(n5310), .D(\vrf/N76 ), .Q(
        \vrf/regTable[1][58] ) );
  LHQD1BWP \vrf/regTable_reg[1][59]  ( .E(n5310), .D(\vrf/N77 ), .Q(
        \vrf/regTable[1][59] ) );
  LHQD1BWP \vrf/regTable_reg[1][60]  ( .E(n5310), .D(\vrf/N78 ), .Q(
        \vrf/regTable[1][60] ) );
  LHQD1BWP \vrf/regTable_reg[1][61]  ( .E(n5310), .D(\vrf/N79 ), .Q(
        \vrf/regTable[1][61] ) );
  LHQD1BWP \vrf/regTable_reg[1][62]  ( .E(n5310), .D(\vrf/N80 ), .Q(
        \vrf/regTable[1][62] ) );
  LHQD1BWP \vrf/regTable_reg[1][63]  ( .E(n5310), .D(\vrf/N81 ), .Q(
        \vrf/regTable[1][63] ) );
  LHQD1BWP \vrf/regTable_reg[1][64]  ( .E(n5310), .D(\vrf/N82 ), .Q(
        \vrf/regTable[1][64] ) );
  LHQD1BWP \vrf/regTable_reg[1][65]  ( .E(n5310), .D(\vrf/N83 ), .Q(
        \vrf/regTable[1][65] ) );
  LHQD1BWP \vrf/regTable_reg[1][66]  ( .E(n5310), .D(\vrf/N84 ), .Q(
        \vrf/regTable[1][66] ) );
  LHQD1BWP \vrf/regTable_reg[1][67]  ( .E(n5310), .D(\vrf/N85 ), .Q(
        \vrf/regTable[1][67] ) );
  LHQD1BWP \vrf/regTable_reg[1][68]  ( .E(n5309), .D(\vrf/N86 ), .Q(
        \vrf/regTable[1][68] ) );
  LHQD1BWP \vrf/regTable_reg[1][69]  ( .E(n5309), .D(\vrf/N87 ), .Q(
        \vrf/regTable[1][69] ) );
  LHQD1BWP \vrf/regTable_reg[1][70]  ( .E(n5309), .D(\vrf/N88 ), .Q(
        \vrf/regTable[1][70] ) );
  LHQD1BWP \vrf/regTable_reg[1][71]  ( .E(n5309), .D(\vrf/N89 ), .Q(
        \vrf/regTable[1][71] ) );
  LHQD1BWP \vrf/regTable_reg[1][72]  ( .E(n5309), .D(\vrf/N90 ), .Q(
        \vrf/regTable[1][72] ) );
  LHQD1BWP \vrf/regTable_reg[1][73]  ( .E(n5309), .D(\vrf/N91 ), .Q(
        \vrf/regTable[1][73] ) );
  LHQD1BWP \vrf/regTable_reg[1][74]  ( .E(n5309), .D(\vrf/N92 ), .Q(
        \vrf/regTable[1][74] ) );
  LHQD1BWP \vrf/regTable_reg[1][75]  ( .E(n5309), .D(\vrf/N93 ), .Q(
        \vrf/regTable[1][75] ) );
  LHQD1BWP \vrf/regTable_reg[1][76]  ( .E(n5309), .D(\vrf/N94 ), .Q(
        \vrf/regTable[1][76] ) );
  LHQD1BWP \vrf/regTable_reg[1][77]  ( .E(n5309), .D(\vrf/N95 ), .Q(
        \vrf/regTable[1][77] ) );
  LHQD1BWP \vrf/regTable_reg[1][78]  ( .E(n5309), .D(\vrf/N96 ), .Q(
        \vrf/regTable[1][78] ) );
  LHQD1BWP \vrf/regTable_reg[1][79]  ( .E(n5308), .D(\vrf/N97 ), .Q(
        \vrf/regTable[1][79] ) );
  LHQD1BWP \vrf/regTable_reg[1][80]  ( .E(n5308), .D(\vrf/N98 ), .Q(
        \vrf/regTable[1][80] ) );
  LHQD1BWP \vrf/regTable_reg[1][81]  ( .E(n5308), .D(\vrf/N99 ), .Q(
        \vrf/regTable[1][81] ) );
  LHQD1BWP \vrf/regTable_reg[1][82]  ( .E(n5308), .D(\vrf/N100 ), .Q(
        \vrf/regTable[1][82] ) );
  LHQD1BWP \vrf/regTable_reg[1][83]  ( .E(n5308), .D(\vrf/N101 ), .Q(
        \vrf/regTable[1][83] ) );
  LHQD1BWP \vrf/regTable_reg[1][84]  ( .E(n5308), .D(\vrf/N102 ), .Q(
        \vrf/regTable[1][84] ) );
  LHQD1BWP \vrf/regTable_reg[1][85]  ( .E(n5308), .D(\vrf/N103 ), .Q(
        \vrf/regTable[1][85] ) );
  LHQD1BWP \vrf/regTable_reg[1][86]  ( .E(n5308), .D(\vrf/N104 ), .Q(
        \vrf/regTable[1][86] ) );
  LHQD1BWP \vrf/regTable_reg[1][87]  ( .E(n5308), .D(\vrf/N105 ), .Q(
        \vrf/regTable[1][87] ) );
  LHQD1BWP \vrf/regTable_reg[1][88]  ( .E(n5308), .D(\vrf/N106 ), .Q(
        \vrf/regTable[1][88] ) );
  LHQD1BWP \vrf/regTable_reg[1][89]  ( .E(n5308), .D(\vrf/N107 ), .Q(
        \vrf/regTable[1][89] ) );
  LHQD1BWP \vrf/regTable_reg[1][90]  ( .E(n5307), .D(\vrf/N108 ), .Q(
        \vrf/regTable[1][90] ) );
  LHQD1BWP \vrf/regTable_reg[1][91]  ( .E(n5307), .D(\vrf/N109 ), .Q(
        \vrf/regTable[1][91] ) );
  LHQD1BWP \vrf/regTable_reg[1][92]  ( .E(n5307), .D(\vrf/N110 ), .Q(
        \vrf/regTable[1][92] ) );
  LHQD1BWP \vrf/regTable_reg[1][93]  ( .E(n5307), .D(\vrf/N111 ), .Q(
        \vrf/regTable[1][93] ) );
  LHQD1BWP \vrf/regTable_reg[1][94]  ( .E(n5307), .D(\vrf/N112 ), .Q(
        \vrf/regTable[1][94] ) );
  LHQD1BWP \vrf/regTable_reg[1][95]  ( .E(n5307), .D(\vrf/N113 ), .Q(
        \vrf/regTable[1][95] ) );
  LHQD1BWP \vrf/regTable_reg[1][96]  ( .E(n5307), .D(\vrf/N114 ), .Q(
        \vrf/regTable[1][96] ) );
  LHQD1BWP \vrf/regTable_reg[1][97]  ( .E(n5307), .D(\vrf/N115 ), .Q(
        \vrf/regTable[1][97] ) );
  LHQD1BWP \vrf/regTable_reg[1][98]  ( .E(n5307), .D(\vrf/N116 ), .Q(
        \vrf/regTable[1][98] ) );
  LHQD1BWP \vrf/regTable_reg[1][99]  ( .E(n5307), .D(\vrf/N118 ), .Q(
        \vrf/regTable[1][99] ) );
  LHQD1BWP \vrf/regTable_reg[1][100]  ( .E(n5317), .D(\vrf/N119 ), .Q(
        \vrf/regTable[1][100] ) );
  LHQD1BWP \vrf/regTable_reg[1][101]  ( .E(n5317), .D(\vrf/N120 ), .Q(
        \vrf/regTable[1][101] ) );
  LHQD1BWP \vrf/regTable_reg[1][102]  ( .E(n5317), .D(\vrf/N121 ), .Q(
        \vrf/regTable[1][102] ) );
  LHQD1BWP \vrf/regTable_reg[1][103]  ( .E(n5317), .D(\vrf/N122 ), .Q(
        \vrf/regTable[1][103] ) );
  LHQD1BWP \vrf/regTable_reg[1][104]  ( .E(n5317), .D(\vrf/N123 ), .Q(
        \vrf/regTable[1][104] ) );
  LHQD1BWP \vrf/regTable_reg[1][105]  ( .E(n5316), .D(\vrf/N124 ), .Q(
        \vrf/regTable[1][105] ) );
  LHQD1BWP \vrf/regTable_reg[1][106]  ( .E(n5316), .D(\vrf/N125 ), .Q(
        \vrf/regTable[1][106] ) );
  LHQD1BWP \vrf/regTable_reg[1][107]  ( .E(n5316), .D(\vrf/N126 ), .Q(
        \vrf/regTable[1][107] ) );
  LHQD1BWP \vrf/regTable_reg[1][108]  ( .E(n5316), .D(\vrf/N127 ), .Q(
        \vrf/regTable[1][108] ) );
  LHQD1BWP \vrf/regTable_reg[1][109]  ( .E(n5316), .D(\vrf/N128 ), .Q(
        \vrf/regTable[1][109] ) );
  LHQD1BWP \vrf/regTable_reg[1][110]  ( .E(n5316), .D(\vrf/N129 ), .Q(
        \vrf/regTable[1][110] ) );
  LHQD1BWP \vrf/regTable_reg[1][111]  ( .E(n5316), .D(\vrf/N130 ), .Q(
        \vrf/regTable[1][111] ) );
  LHQD1BWP \vrf/regTable_reg[1][112]  ( .E(n5316), .D(\vrf/N131 ), .Q(
        \vrf/regTable[1][112] ) );
  LHQD1BWP \vrf/regTable_reg[1][113]  ( .E(n5316), .D(\vrf/N132 ), .Q(
        \vrf/regTable[1][113] ) );
  LHQD1BWP \vrf/regTable_reg[1][114]  ( .E(n5316), .D(\vrf/N133 ), .Q(
        \vrf/regTable[1][114] ) );
  LHQD1BWP \vrf/regTable_reg[1][115]  ( .E(n5316), .D(\vrf/N134 ), .Q(
        \vrf/regTable[1][115] ) );
  LHQD1BWP \vrf/regTable_reg[1][116]  ( .E(n5315), .D(\vrf/N135 ), .Q(
        \vrf/regTable[1][116] ) );
  LHQD1BWP \vrf/regTable_reg[1][117]  ( .E(n5315), .D(\vrf/N136 ), .Q(
        \vrf/regTable[1][117] ) );
  LHQD1BWP \vrf/regTable_reg[1][118]  ( .E(n5315), .D(\vrf/N137 ), .Q(
        \vrf/regTable[1][118] ) );
  LHQD1BWP \vrf/regTable_reg[1][119]  ( .E(n5315), .D(\vrf/N138 ), .Q(
        \vrf/regTable[1][119] ) );
  LHQD1BWP \vrf/regTable_reg[1][120]  ( .E(n5315), .D(\vrf/N139 ), .Q(
        \vrf/regTable[1][120] ) );
  LHQD1BWP \vrf/regTable_reg[1][121]  ( .E(n5315), .D(\vrf/N140 ), .Q(
        \vrf/regTable[1][121] ) );
  LHQD1BWP \vrf/regTable_reg[1][122]  ( .E(n5315), .D(\vrf/N141 ), .Q(
        \vrf/regTable[1][122] ) );
  LHQD1BWP \vrf/regTable_reg[1][123]  ( .E(n5315), .D(\vrf/N142 ), .Q(
        \vrf/regTable[1][123] ) );
  LHQD1BWP \vrf/regTable_reg[1][124]  ( .E(n5315), .D(\vrf/N143 ), .Q(
        \vrf/regTable[1][124] ) );
  LHQD1BWP \vrf/regTable_reg[1][125]  ( .E(n5315), .D(\vrf/N144 ), .Q(
        \vrf/regTable[1][125] ) );
  LHQD1BWP \vrf/regTable_reg[1][126]  ( .E(n5315), .D(\vrf/N145 ), .Q(
        \vrf/regTable[1][126] ) );
  LHQD1BWP \vrf/regTable_reg[1][127]  ( .E(n5314), .D(\vrf/N146 ), .Q(
        \vrf/regTable[1][127] ) );
  LHQD1BWP \vrf/regTable_reg[1][128]  ( .E(n5317), .D(\vrf/N147 ), .Q(
        \vrf/regTable[1][128] ) );
  LHQD1BWP \vrf/regTable_reg[1][129]  ( .E(n5317), .D(\vrf/N148 ), .Q(
        \vrf/regTable[1][129] ) );
  LHQD1BWP \vrf/regTable_reg[1][130]  ( .E(n5317), .D(\vrf/N149 ), .Q(
        \vrf/regTable[1][130] ) );
  LHQD1BWP \vrf/regTable_reg[1][131]  ( .E(n5317), .D(\vrf/N150 ), .Q(
        \vrf/regTable[1][131] ) );
  LHQD1BWP \vrf/regTable_reg[1][132]  ( .E(n5317), .D(\vrf/N151 ), .Q(
        \vrf/regTable[1][132] ) );
  LHQD1BWP \vrf/regTable_reg[1][133]  ( .E(n5317), .D(\vrf/N152 ), .Q(
        \vrf/regTable[1][133] ) );
  LHQD1BWP \vrf/regTable_reg[1][134]  ( .E(n5318), .D(\vrf/N153 ), .Q(
        \vrf/regTable[1][134] ) );
  LHQD1BWP \vrf/regTable_reg[1][135]  ( .E(n5318), .D(\vrf/N154 ), .Q(
        \vrf/regTable[1][135] ) );
  LHQD1BWP \vrf/regTable_reg[1][136]  ( .E(n5318), .D(\vrf/N155 ), .Q(
        \vrf/regTable[1][136] ) );
  LHQD1BWP \vrf/regTable_reg[1][137]  ( .E(n5318), .D(\vrf/N156 ), .Q(
        \vrf/regTable[1][137] ) );
  LHQD1BWP \vrf/regTable_reg[1][138]  ( .E(n5318), .D(\vrf/N157 ), .Q(
        \vrf/regTable[1][138] ) );
  LHQD1BWP \vrf/regTable_reg[1][139]  ( .E(n5318), .D(\vrf/N158 ), .Q(
        \vrf/regTable[1][139] ) );
  LHQD1BWP \vrf/regTable_reg[1][140]  ( .E(n5318), .D(\vrf/N159 ), .Q(
        \vrf/regTable[1][140] ) );
  LHQD1BWP \vrf/regTable_reg[1][141]  ( .E(n5318), .D(\vrf/N160 ), .Q(
        \vrf/regTable[1][141] ) );
  LHQD1BWP \vrf/regTable_reg[1][142]  ( .E(n5318), .D(\vrf/N161 ), .Q(
        \vrf/regTable[1][142] ) );
  LHQD1BWP \vrf/regTable_reg[1][143]  ( .E(n5318), .D(\vrf/N162 ), .Q(
        \vrf/regTable[1][143] ) );
  LHQD1BWP \vrf/regTable_reg[1][144]  ( .E(n5318), .D(\vrf/N163 ), .Q(
        \vrf/regTable[1][144] ) );
  LHQD1BWP \vrf/regTable_reg[1][145]  ( .E(n5318), .D(\vrf/N164 ), .Q(
        \vrf/regTable[1][145] ) );
  LHQD1BWP \vrf/regTable_reg[1][146]  ( .E(n5319), .D(\vrf/N165 ), .Q(
        \vrf/regTable[1][146] ) );
  LHQD1BWP \vrf/regTable_reg[1][147]  ( .E(n5319), .D(\vrf/N166 ), .Q(
        \vrf/regTable[1][147] ) );
  LHQD1BWP \vrf/regTable_reg[1][148]  ( .E(n5319), .D(\vrf/N167 ), .Q(
        \vrf/regTable[1][148] ) );
  LHQD1BWP \vrf/regTable_reg[1][149]  ( .E(n5319), .D(\vrf/N168 ), .Q(
        \vrf/regTable[1][149] ) );
  LHQD1BWP \vrf/regTable_reg[1][150]  ( .E(n5319), .D(\vrf/N169 ), .Q(
        \vrf/regTable[1][150] ) );
  LHQD1BWP \vrf/regTable_reg[1][151]  ( .E(n5319), .D(\vrf/N170 ), .Q(
        \vrf/regTable[1][151] ) );
  LHQD1BWP \vrf/regTable_reg[1][152]  ( .E(n5319), .D(\vrf/N171 ), .Q(
        \vrf/regTable[1][152] ) );
  LHQD1BWP \vrf/regTable_reg[1][153]  ( .E(n5319), .D(\vrf/N172 ), .Q(
        \vrf/regTable[1][153] ) );
  LHQD1BWP \vrf/regTable_reg[1][154]  ( .E(n5319), .D(\vrf/N173 ), .Q(
        \vrf/regTable[1][154] ) );
  LHQD1BWP \vrf/regTable_reg[1][155]  ( .E(n5319), .D(\vrf/N174 ), .Q(
        \vrf/regTable[1][155] ) );
  LHQD1BWP \vrf/regTable_reg[1][156]  ( .E(n5319), .D(\vrf/N175 ), .Q(
        \vrf/regTable[1][156] ) );
  LHQD1BWP \vrf/regTable_reg[1][157]  ( .E(n5319), .D(\vrf/N176 ), .Q(
        \vrf/regTable[1][157] ) );
  LHQD1BWP \vrf/regTable_reg[1][158]  ( .E(n5320), .D(\vrf/N177 ), .Q(
        \vrf/regTable[1][158] ) );
  LHQD1BWP \vrf/regTable_reg[1][159]  ( .E(n5320), .D(\vrf/N178 ), .Q(
        \vrf/regTable[1][159] ) );
  LHQD1BWP \vrf/regTable_reg[1][160]  ( .E(n5320), .D(\vrf/N179 ), .Q(
        \vrf/regTable[1][160] ) );
  LHQD1BWP \vrf/regTable_reg[1][161]  ( .E(n5320), .D(\vrf/N180 ), .Q(
        \vrf/regTable[1][161] ) );
  LHQD1BWP \vrf/regTable_reg[1][162]  ( .E(n5320), .D(\vrf/N181 ), .Q(
        \vrf/regTable[1][162] ) );
  LHQD1BWP \vrf/regTable_reg[1][163]  ( .E(n5320), .D(\vrf/N182 ), .Q(
        \vrf/regTable[1][163] ) );
  LHQD1BWP \vrf/regTable_reg[1][164]  ( .E(n5320), .D(\vrf/N183 ), .Q(
        \vrf/regTable[1][164] ) );
  LHQD1BWP \vrf/regTable_reg[1][165]  ( .E(n5320), .D(\vrf/N184 ), .Q(
        \vrf/regTable[1][165] ) );
  LHQD1BWP \vrf/regTable_reg[1][166]  ( .E(n5320), .D(\vrf/N185 ), .Q(
        \vrf/regTable[1][166] ) );
  LHQD1BWP \vrf/regTable_reg[1][167]  ( .E(n5320), .D(\vrf/N186 ), .Q(
        \vrf/regTable[1][167] ) );
  LHQD1BWP \vrf/regTable_reg[1][168]  ( .E(n5320), .D(\vrf/N187 ), .Q(
        \vrf/regTable[1][168] ) );
  LHQD1BWP \vrf/regTable_reg[1][169]  ( .E(n5320), .D(\vrf/N188 ), .Q(
        \vrf/regTable[1][169] ) );
  LHQD1BWP \vrf/regTable_reg[1][170]  ( .E(n5321), .D(\vrf/N189 ), .Q(
        \vrf/regTable[1][170] ) );
  LHQD1BWP \vrf/regTable_reg[1][171]  ( .E(n5321), .D(\vrf/N190 ), .Q(
        \vrf/regTable[1][171] ) );
  LHQD1BWP \vrf/regTable_reg[1][172]  ( .E(n5321), .D(\vrf/N191 ), .Q(
        \vrf/regTable[1][172] ) );
  LHQD1BWP \vrf/regTable_reg[1][173]  ( .E(n5321), .D(\vrf/N192 ), .Q(
        \vrf/regTable[1][173] ) );
  LHQD1BWP \vrf/regTable_reg[1][174]  ( .E(n5321), .D(\vrf/N193 ), .Q(
        \vrf/regTable[1][174] ) );
  LHQD1BWP \vrf/regTable_reg[1][175]  ( .E(n5321), .D(\vrf/N194 ), .Q(
        \vrf/regTable[1][175] ) );
  LHQD1BWP \vrf/regTable_reg[1][176]  ( .E(n5321), .D(\vrf/N195 ), .Q(
        \vrf/regTable[1][176] ) );
  LHQD1BWP \vrf/regTable_reg[1][177]  ( .E(n5321), .D(\vrf/N196 ), .Q(
        \vrf/regTable[1][177] ) );
  LHQD1BWP \vrf/regTable_reg[1][178]  ( .E(n5321), .D(\vrf/N197 ), .Q(
        \vrf/regTable[1][178] ) );
  LHQD1BWP \vrf/regTable_reg[1][179]  ( .E(n5321), .D(\vrf/N198 ), .Q(
        \vrf/regTable[1][179] ) );
  LHQD1BWP \vrf/regTable_reg[1][180]  ( .E(n5321), .D(\vrf/N199 ), .Q(
        \vrf/regTable[1][180] ) );
  LHQD1BWP \vrf/regTable_reg[1][181]  ( .E(n5321), .D(\vrf/N200 ), .Q(
        \vrf/regTable[1][181] ) );
  LHQD1BWP \vrf/regTable_reg[1][182]  ( .E(n5322), .D(\vrf/N201 ), .Q(
        \vrf/regTable[1][182] ) );
  LHQD1BWP \vrf/regTable_reg[1][183]  ( .E(n5322), .D(\vrf/N202 ), .Q(
        \vrf/regTable[1][183] ) );
  LHQD1BWP \vrf/regTable_reg[1][184]  ( .E(n5322), .D(\vrf/N203 ), .Q(
        \vrf/regTable[1][184] ) );
  LHQD1BWP \vrf/regTable_reg[1][185]  ( .E(n5322), .D(\vrf/N204 ), .Q(
        \vrf/regTable[1][185] ) );
  LHQD1BWP \vrf/regTable_reg[1][186]  ( .E(n5322), .D(\vrf/N205 ), .Q(
        \vrf/regTable[1][186] ) );
  LHQD1BWP \vrf/regTable_reg[1][187]  ( .E(n5322), .D(\vrf/N206 ), .Q(
        \vrf/regTable[1][187] ) );
  LHQD1BWP \vrf/regTable_reg[1][188]  ( .E(n5322), .D(\vrf/N207 ), .Q(
        \vrf/regTable[1][188] ) );
  LHQD1BWP \vrf/regTable_reg[1][189]  ( .E(n5322), .D(\vrf/N208 ), .Q(
        \vrf/regTable[1][189] ) );
  LHQD1BWP \vrf/regTable_reg[1][190]  ( .E(n5322), .D(\vrf/N209 ), .Q(
        \vrf/regTable[1][190] ) );
  LHQD1BWP \vrf/regTable_reg[1][191]  ( .E(n5322), .D(\vrf/N210 ), .Q(
        \vrf/regTable[1][191] ) );
  LHQD1BWP \vrf/regTable_reg[1][192]  ( .E(n5322), .D(\vrf/N211 ), .Q(
        \vrf/regTable[1][192] ) );
  LHQD1BWP \vrf/regTable_reg[1][193]  ( .E(n5322), .D(\vrf/N212 ), .Q(
        \vrf/regTable[1][193] ) );
  LHQD1BWP \vrf/regTable_reg[1][194]  ( .E(n5323), .D(\vrf/N213 ), .Q(
        \vrf/regTable[1][194] ) );
  LHQD1BWP \vrf/regTable_reg[1][195]  ( .E(n5323), .D(\vrf/N214 ), .Q(
        \vrf/regTable[1][195] ) );
  LHQD1BWP \vrf/regTable_reg[1][196]  ( .E(n5323), .D(\vrf/N215 ), .Q(
        \vrf/regTable[1][196] ) );
  LHQD1BWP \vrf/regTable_reg[1][197]  ( .E(n5323), .D(\vrf/N216 ), .Q(
        \vrf/regTable[1][197] ) );
  LHQD1BWP \vrf/regTable_reg[1][198]  ( .E(n5323), .D(\vrf/N218 ), .Q(
        \vrf/regTable[1][198] ) );
  LHQD1BWP \vrf/regTable_reg[1][199]  ( .E(n5323), .D(\vrf/N219 ), .Q(
        \vrf/regTable[1][199] ) );
  LHQD1BWP \vrf/regTable_reg[1][200]  ( .E(n5323), .D(\vrf/N220 ), .Q(
        \vrf/regTable[1][200] ) );
  LHQD1BWP \vrf/regTable_reg[1][201]  ( .E(n5323), .D(\vrf/N221 ), .Q(
        \vrf/regTable[1][201] ) );
  LHQD1BWP \vrf/regTable_reg[1][202]  ( .E(n5323), .D(\vrf/N222 ), .Q(
        \vrf/regTable[1][202] ) );
  LHQD1BWP \vrf/regTable_reg[1][203]  ( .E(n5323), .D(\vrf/N223 ), .Q(
        \vrf/regTable[1][203] ) );
  LHQD1BWP \vrf/regTable_reg[1][204]  ( .E(n5323), .D(\vrf/N224 ), .Q(
        \vrf/regTable[1][204] ) );
  LHQD1BWP \vrf/regTable_reg[1][205]  ( .E(n5323), .D(\vrf/N225 ), .Q(
        \vrf/regTable[1][205] ) );
  LHQD1BWP \vrf/regTable_reg[1][206]  ( .E(n5324), .D(\vrf/N226 ), .Q(
        \vrf/regTable[1][206] ) );
  LHQD1BWP \vrf/regTable_reg[1][207]  ( .E(n5324), .D(\vrf/N227 ), .Q(
        \vrf/regTable[1][207] ) );
  LHQD1BWP \vrf/regTable_reg[1][208]  ( .E(n5324), .D(\vrf/N228 ), .Q(
        \vrf/regTable[1][208] ) );
  LHQD1BWP \vrf/regTable_reg[1][209]  ( .E(n5324), .D(\vrf/N229 ), .Q(
        \vrf/regTable[1][209] ) );
  LHQD1BWP \vrf/regTable_reg[1][210]  ( .E(n5324), .D(\vrf/N230 ), .Q(
        \vrf/regTable[1][210] ) );
  LHQD1BWP \vrf/regTable_reg[1][211]  ( .E(n5324), .D(\vrf/N231 ), .Q(
        \vrf/regTable[1][211] ) );
  LHQD1BWP \vrf/regTable_reg[1][212]  ( .E(n5324), .D(\vrf/N232 ), .Q(
        \vrf/regTable[1][212] ) );
  LHQD1BWP \vrf/regTable_reg[1][213]  ( .E(n5324), .D(\vrf/N233 ), .Q(
        \vrf/regTable[1][213] ) );
  LHQD1BWP \vrf/regTable_reg[1][214]  ( .E(n5324), .D(\vrf/N234 ), .Q(
        \vrf/regTable[1][214] ) );
  LHQD1BWP \vrf/regTable_reg[1][215]  ( .E(n5324), .D(\vrf/N235 ), .Q(
        \vrf/regTable[1][215] ) );
  LHQD1BWP \vrf/regTable_reg[1][216]  ( .E(n5324), .D(\vrf/N236 ), .Q(
        \vrf/regTable[1][216] ) );
  LHQD1BWP \vrf/regTable_reg[1][217]  ( .E(n5324), .D(\vrf/N237 ), .Q(
        \vrf/regTable[1][217] ) );
  LHQD1BWP \vrf/regTable_reg[1][218]  ( .E(n5325), .D(\vrf/N238 ), .Q(
        \vrf/regTable[1][218] ) );
  LHQD1BWP \vrf/regTable_reg[1][219]  ( .E(n5325), .D(\vrf/N239 ), .Q(
        \vrf/regTable[1][219] ) );
  LHQD1BWP \vrf/regTable_reg[1][220]  ( .E(n5325), .D(\vrf/N240 ), .Q(
        \vrf/regTable[1][220] ) );
  LHQD1BWP \vrf/regTable_reg[1][221]  ( .E(n5325), .D(\vrf/N241 ), .Q(
        \vrf/regTable[1][221] ) );
  LHQD1BWP \vrf/regTable_reg[1][222]  ( .E(n5325), .D(\vrf/N242 ), .Q(
        \vrf/regTable[1][222] ) );
  LHQD1BWP \vrf/regTable_reg[1][223]  ( .E(n5325), .D(\vrf/N243 ), .Q(
        \vrf/regTable[1][223] ) );
  LHQD1BWP \vrf/regTable_reg[1][224]  ( .E(n5325), .D(\vrf/N244 ), .Q(
        \vrf/regTable[1][224] ) );
  LHQD1BWP \vrf/regTable_reg[1][225]  ( .E(n5325), .D(\vrf/N245 ), .Q(
        \vrf/regTable[1][225] ) );
  LHQD1BWP \vrf/regTable_reg[1][226]  ( .E(n5325), .D(\vrf/N246 ), .Q(
        \vrf/regTable[1][226] ) );
  LHQD1BWP \vrf/regTable_reg[1][227]  ( .E(n5325), .D(\vrf/N247 ), .Q(
        \vrf/regTable[1][227] ) );
  LHQD1BWP \vrf/regTable_reg[1][228]  ( .E(n5325), .D(\vrf/N248 ), .Q(
        \vrf/regTable[1][228] ) );
  LHQD1BWP \vrf/regTable_reg[1][229]  ( .E(n5325), .D(\vrf/N249 ), .Q(
        \vrf/regTable[1][229] ) );
  LHQD1BWP \vrf/regTable_reg[1][230]  ( .E(n5326), .D(\vrf/N250 ), .Q(
        \vrf/regTable[1][230] ) );
  LHQD1BWP \vrf/regTable_reg[1][231]  ( .E(n5326), .D(\vrf/N251 ), .Q(
        \vrf/regTable[1][231] ) );
  LHQD1BWP \vrf/regTable_reg[1][232]  ( .E(n5326), .D(\vrf/N252 ), .Q(
        \vrf/regTable[1][232] ) );
  LHQD1BWP \vrf/regTable_reg[1][233]  ( .E(n5326), .D(\vrf/N253 ), .Q(
        \vrf/regTable[1][233] ) );
  LHQD1BWP \vrf/regTable_reg[1][234]  ( .E(n5326), .D(\vrf/N254 ), .Q(
        \vrf/regTable[1][234] ) );
  LHQD1BWP \vrf/regTable_reg[1][235]  ( .E(n5326), .D(\vrf/N255 ), .Q(
        \vrf/regTable[1][235] ) );
  LHQD1BWP \vrf/regTable_reg[1][236]  ( .E(n5326), .D(\vrf/N256 ), .Q(
        \vrf/regTable[1][236] ) );
  LHQD1BWP \vrf/regTable_reg[1][237]  ( .E(n5326), .D(\vrf/N257 ), .Q(
        \vrf/regTable[1][237] ) );
  LHQD1BWP \vrf/regTable_reg[1][238]  ( .E(n5326), .D(\vrf/N258 ), .Q(
        \vrf/regTable[1][238] ) );
  LHQD1BWP \vrf/regTable_reg[1][239]  ( .E(n5326), .D(\vrf/N259 ), .Q(
        \vrf/regTable[1][239] ) );
  LHQD1BWP \vrf/regTable_reg[1][240]  ( .E(n5326), .D(\vrf/N260 ), .Q(
        \vrf/regTable[1][240] ) );
  LHQD1BWP \vrf/regTable_reg[1][241]  ( .E(n5326), .D(\vrf/N261 ), .Q(
        \vrf/regTable[1][241] ) );
  LHQD1BWP \vrf/regTable_reg[1][242]  ( .E(n5327), .D(\vrf/N262 ), .Q(
        \vrf/regTable[1][242] ) );
  LHQD1BWP \vrf/regTable_reg[1][243]  ( .E(n5327), .D(\vrf/N263 ), .Q(
        \vrf/regTable[1][243] ) );
  LHQD1BWP \vrf/regTable_reg[1][244]  ( .E(n5327), .D(\vrf/N264 ), .Q(
        \vrf/regTable[1][244] ) );
  LHQD1BWP \vrf/regTable_reg[1][245]  ( .E(n5327), .D(\vrf/N265 ), .Q(
        \vrf/regTable[1][245] ) );
  LHQD1BWP \vrf/regTable_reg[1][246]  ( .E(n5327), .D(\vrf/N266 ), .Q(
        \vrf/regTable[1][246] ) );
  LHQD1BWP \vrf/regTable_reg[1][247]  ( .E(n5327), .D(\vrf/N267 ), .Q(
        \vrf/regTable[1][247] ) );
  LHQD1BWP \vrf/regTable_reg[1][248]  ( .E(n5327), .D(\vrf/N268 ), .Q(
        \vrf/regTable[1][248] ) );
  LHQD1BWP \vrf/regTable_reg[1][249]  ( .E(n5327), .D(\vrf/N269 ), .Q(
        \vrf/regTable[1][249] ) );
  LHQD1BWP \vrf/regTable_reg[1][250]  ( .E(n5327), .D(\vrf/N270 ), .Q(
        \vrf/regTable[1][250] ) );
  LHQD1BWP \vrf/regTable_reg[1][251]  ( .E(n5327), .D(\vrf/N271 ), .Q(
        \vrf/regTable[1][251] ) );
  LHQD1BWP \vrf/regTable_reg[1][252]  ( .E(n5327), .D(\vrf/N272 ), .Q(
        \vrf/regTable[1][252] ) );
  LHQD1BWP \vrf/regTable_reg[1][253]  ( .E(n5327), .D(\vrf/N273 ), .Q(
        \vrf/regTable[1][253] ) );
  LHQD1BWP \vrf/regTable_reg[6][15]  ( .E(n5158), .D(\vrf/N33 ), .Q(
        \vrf/regTable[6][15] ) );
  LHQD1BWP \vrf/regTable_reg[6][16]  ( .E(n5158), .D(\vrf/N34 ), .Q(
        \vrf/regTable[6][16] ) );
  LHQD1BWP \vrf/regTable_reg[6][254]  ( .E(n5158), .D(\vrf/N274 ), .Q(
        \vrf/regTable[6][254] ) );
  LHQD1BWP \vrf/regTable_reg[6][255]  ( .E(n5158), .D(\vrf/N275 ), .Q(
        \vrf/regTable[6][255] ) );
  LHQD1BWP \vrf/regTable_reg[2][15]  ( .E(n5294), .D(\vrf/N33 ), .Q(
        \vrf/regTable[2][15] ) );
  LHQD1BWP \vrf/regTable_reg[2][16]  ( .E(n5294), .D(\vrf/N34 ), .Q(
        \vrf/regTable[2][16] ) );
  LHQD1BWP \vrf/regTable_reg[2][254]  ( .E(n5294), .D(\vrf/N274 ), .Q(
        \vrf/regTable[2][254] ) );
  LHQD1BWP \vrf/regTable_reg[2][255]  ( .E(n5294), .D(\vrf/N275 ), .Q(
        \vrf/regTable[2][255] ) );
  LHQD1BWP \vrf/regTable_reg[6][0]  ( .E(n5147), .D(\vrf/N18 ), .Q(
        \vrf/regTable[6][0] ) );
  LHQD1BWP \vrf/regTable_reg[6][1]  ( .E(n5144), .D(\vrf/N19 ), .Q(
        \vrf/regTable[6][1] ) );
  LHQD1BWP \vrf/regTable_reg[6][2]  ( .E(n5143), .D(\vrf/N20 ), .Q(
        \vrf/regTable[6][2] ) );
  LHQD1BWP \vrf/regTable_reg[6][3]  ( .E(n5142), .D(\vrf/N21 ), .Q(
        \vrf/regTable[6][3] ) );
  LHQD1BWP \vrf/regTable_reg[6][4]  ( .E(n5141), .D(\vrf/N22 ), .Q(
        \vrf/regTable[6][4] ) );
  LHQD1BWP \vrf/regTable_reg[6][5]  ( .E(n5140), .D(\vrf/N23 ), .Q(
        \vrf/regTable[6][5] ) );
  LHQD1BWP \vrf/regTable_reg[6][6]  ( .E(n5139), .D(\vrf/N24 ), .Q(
        \vrf/regTable[6][6] ) );
  LHQD1BWP \vrf/regTable_reg[6][7]  ( .E(n5138), .D(\vrf/N25 ), .Q(
        \vrf/regTable[6][7] ) );
  LHQD1BWP \vrf/regTable_reg[6][8]  ( .E(n5137), .D(\vrf/N26 ), .Q(
        \vrf/regTable[6][8] ) );
  LHQD1BWP \vrf/regTable_reg[6][9]  ( .E(n5137), .D(\vrf/N27 ), .Q(
        \vrf/regTable[6][9] ) );
  LHQD1BWP \vrf/regTable_reg[6][10]  ( .E(n5146), .D(\vrf/N28 ), .Q(
        \vrf/regTable[6][10] ) );
  LHQD1BWP \vrf/regTable_reg[6][11]  ( .E(n5145), .D(\vrf/N29 ), .Q(
        \vrf/regTable[6][11] ) );
  LHQD1BWP \vrf/regTable_reg[6][12]  ( .E(n5144), .D(\vrf/N30 ), .Q(
        \vrf/regTable[6][12] ) );
  LHQD1BWP \vrf/regTable_reg[6][13]  ( .E(n5144), .D(\vrf/N31 ), .Q(
        \vrf/regTable[6][13] ) );
  LHQD1BWP \vrf/regTable_reg[6][14]  ( .E(n5144), .D(\vrf/N32 ), .Q(
        \vrf/regTable[6][14] ) );
  LHQD1BWP \vrf/regTable_reg[6][17]  ( .E(n5144), .D(\vrf/N35 ), .Q(
        \vrf/regTable[6][17] ) );
  LHQD1BWP \vrf/regTable_reg[6][18]  ( .E(n5144), .D(\vrf/N36 ), .Q(
        \vrf/regTable[6][18] ) );
  LHQD1BWP \vrf/regTable_reg[6][19]  ( .E(n5144), .D(\vrf/N37 ), .Q(
        \vrf/regTable[6][19] ) );
  LHQD1BWP \vrf/regTable_reg[6][20]  ( .E(n5144), .D(\vrf/N38 ), .Q(
        \vrf/regTable[6][20] ) );
  LHQD1BWP \vrf/regTable_reg[6][21]  ( .E(n5144), .D(\vrf/N39 ), .Q(
        \vrf/regTable[6][21] ) );
  LHQD1BWP \vrf/regTable_reg[6][22]  ( .E(n5144), .D(\vrf/N40 ), .Q(
        \vrf/regTable[6][22] ) );
  LHQD1BWP \vrf/regTable_reg[6][23]  ( .E(n5144), .D(\vrf/N41 ), .Q(
        \vrf/regTable[6][23] ) );
  LHQD1BWP \vrf/regTable_reg[6][24]  ( .E(n5143), .D(\vrf/N42 ), .Q(
        \vrf/regTable[6][24] ) );
  LHQD1BWP \vrf/regTable_reg[6][25]  ( .E(n5143), .D(\vrf/N43 ), .Q(
        \vrf/regTable[6][25] ) );
  LHQD1BWP \vrf/regTable_reg[6][26]  ( .E(n5143), .D(\vrf/N44 ), .Q(
        \vrf/regTable[6][26] ) );
  LHQD1BWP \vrf/regTable_reg[6][27]  ( .E(n5143), .D(\vrf/N45 ), .Q(
        \vrf/regTable[6][27] ) );
  LHQD1BWP \vrf/regTable_reg[6][28]  ( .E(n5143), .D(\vrf/N46 ), .Q(
        \vrf/regTable[6][28] ) );
  LHQD1BWP \vrf/regTable_reg[6][29]  ( .E(n5143), .D(\vrf/N47 ), .Q(
        \vrf/regTable[6][29] ) );
  LHQD1BWP \vrf/regTable_reg[6][30]  ( .E(n5143), .D(\vrf/N48 ), .Q(
        \vrf/regTable[6][30] ) );
  LHQD1BWP \vrf/regTable_reg[6][31]  ( .E(n5143), .D(\vrf/N49 ), .Q(
        \vrf/regTable[6][31] ) );
  LHQD1BWP \vrf/regTable_reg[6][32]  ( .E(n5143), .D(\vrf/N50 ), .Q(
        \vrf/regTable[6][32] ) );
  LHQD1BWP \vrf/regTable_reg[6][33]  ( .E(n5143), .D(\vrf/N51 ), .Q(
        \vrf/regTable[6][33] ) );
  LHQD1BWP \vrf/regTable_reg[6][34]  ( .E(n5143), .D(\vrf/N52 ), .Q(
        \vrf/regTable[6][34] ) );
  LHQD1BWP \vrf/regTable_reg[6][35]  ( .E(n5142), .D(\vrf/N53 ), .Q(
        \vrf/regTable[6][35] ) );
  LHQD1BWP \vrf/regTable_reg[6][36]  ( .E(n5142), .D(\vrf/N54 ), .Q(
        \vrf/regTable[6][36] ) );
  LHQD1BWP \vrf/regTable_reg[6][37]  ( .E(n5142), .D(\vrf/N55 ), .Q(
        \vrf/regTable[6][37] ) );
  LHQD1BWP \vrf/regTable_reg[6][38]  ( .E(n5142), .D(\vrf/N56 ), .Q(
        \vrf/regTable[6][38] ) );
  LHQD1BWP \vrf/regTable_reg[6][39]  ( .E(n5142), .D(\vrf/N57 ), .Q(
        \vrf/regTable[6][39] ) );
  LHQD1BWP \vrf/regTable_reg[6][40]  ( .E(n5142), .D(\vrf/N58 ), .Q(
        \vrf/regTable[6][40] ) );
  LHQD1BWP \vrf/regTable_reg[6][41]  ( .E(n5142), .D(\vrf/N59 ), .Q(
        \vrf/regTable[6][41] ) );
  LHQD1BWP \vrf/regTable_reg[6][42]  ( .E(n5142), .D(\vrf/N60 ), .Q(
        \vrf/regTable[6][42] ) );
  LHQD1BWP \vrf/regTable_reg[6][43]  ( .E(n5142), .D(\vrf/N61 ), .Q(
        \vrf/regTable[6][43] ) );
  LHQD1BWP \vrf/regTable_reg[6][44]  ( .E(n5142), .D(\vrf/N62 ), .Q(
        \vrf/regTable[6][44] ) );
  LHQD1BWP \vrf/regTable_reg[6][45]  ( .E(n5142), .D(\vrf/N63 ), .Q(
        \vrf/regTable[6][45] ) );
  LHQD1BWP \vrf/regTable_reg[6][46]  ( .E(n5141), .D(\vrf/N64 ), .Q(
        \vrf/regTable[6][46] ) );
  LHQD1BWP \vrf/regTable_reg[6][47]  ( .E(n5141), .D(\vrf/N65 ), .Q(
        \vrf/regTable[6][47] ) );
  LHQD1BWP \vrf/regTable_reg[6][48]  ( .E(n5141), .D(\vrf/N66 ), .Q(
        \vrf/regTable[6][48] ) );
  LHQD1BWP \vrf/regTable_reg[6][49]  ( .E(n5141), .D(\vrf/N67 ), .Q(
        \vrf/regTable[6][49] ) );
  LHQD1BWP \vrf/regTable_reg[6][50]  ( .E(n5141), .D(\vrf/N68 ), .Q(
        \vrf/regTable[6][50] ) );
  LHQD1BWP \vrf/regTable_reg[6][51]  ( .E(n5141), .D(\vrf/N69 ), .Q(
        \vrf/regTable[6][51] ) );
  LHQD1BWP \vrf/regTable_reg[6][52]  ( .E(n5141), .D(\vrf/N70 ), .Q(
        \vrf/regTable[6][52] ) );
  LHQD1BWP \vrf/regTable_reg[6][53]  ( .E(n5141), .D(\vrf/N71 ), .Q(
        \vrf/regTable[6][53] ) );
  LHQD1BWP \vrf/regTable_reg[6][54]  ( .E(n5141), .D(\vrf/N72 ), .Q(
        \vrf/regTable[6][54] ) );
  LHQD1BWP \vrf/regTable_reg[6][55]  ( .E(n5141), .D(\vrf/N73 ), .Q(
        \vrf/regTable[6][55] ) );
  LHQD1BWP \vrf/regTable_reg[6][56]  ( .E(n5141), .D(\vrf/N74 ), .Q(
        \vrf/regTable[6][56] ) );
  LHQD1BWP \vrf/regTable_reg[6][57]  ( .E(n5140), .D(\vrf/N75 ), .Q(
        \vrf/regTable[6][57] ) );
  LHQD1BWP \vrf/regTable_reg[6][58]  ( .E(n5140), .D(\vrf/N76 ), .Q(
        \vrf/regTable[6][58] ) );
  LHQD1BWP \vrf/regTable_reg[6][59]  ( .E(n5140), .D(\vrf/N77 ), .Q(
        \vrf/regTable[6][59] ) );
  LHQD1BWP \vrf/regTable_reg[6][60]  ( .E(n5140), .D(\vrf/N78 ), .Q(
        \vrf/regTable[6][60] ) );
  LHQD1BWP \vrf/regTable_reg[6][61]  ( .E(n5140), .D(\vrf/N79 ), .Q(
        \vrf/regTable[6][61] ) );
  LHQD1BWP \vrf/regTable_reg[6][62]  ( .E(n5140), .D(\vrf/N80 ), .Q(
        \vrf/regTable[6][62] ) );
  LHQD1BWP \vrf/regTable_reg[6][63]  ( .E(n5140), .D(\vrf/N81 ), .Q(
        \vrf/regTable[6][63] ) );
  LHQD1BWP \vrf/regTable_reg[6][64]  ( .E(n5140), .D(\vrf/N82 ), .Q(
        \vrf/regTable[6][64] ) );
  LHQD1BWP \vrf/regTable_reg[6][65]  ( .E(n5140), .D(\vrf/N83 ), .Q(
        \vrf/regTable[6][65] ) );
  LHQD1BWP \vrf/regTable_reg[6][66]  ( .E(n5140), .D(\vrf/N84 ), .Q(
        \vrf/regTable[6][66] ) );
  LHQD1BWP \vrf/regTable_reg[6][67]  ( .E(n5140), .D(\vrf/N85 ), .Q(
        \vrf/regTable[6][67] ) );
  LHQD1BWP \vrf/regTable_reg[6][68]  ( .E(n5139), .D(\vrf/N86 ), .Q(
        \vrf/regTable[6][68] ) );
  LHQD1BWP \vrf/regTable_reg[6][69]  ( .E(n5139), .D(\vrf/N87 ), .Q(
        \vrf/regTable[6][69] ) );
  LHQD1BWP \vrf/regTable_reg[6][70]  ( .E(n5139), .D(\vrf/N88 ), .Q(
        \vrf/regTable[6][70] ) );
  LHQD1BWP \vrf/regTable_reg[6][71]  ( .E(n5139), .D(\vrf/N89 ), .Q(
        \vrf/regTable[6][71] ) );
  LHQD1BWP \vrf/regTable_reg[6][72]  ( .E(n5139), .D(\vrf/N90 ), .Q(
        \vrf/regTable[6][72] ) );
  LHQD1BWP \vrf/regTable_reg[6][73]  ( .E(n5139), .D(\vrf/N91 ), .Q(
        \vrf/regTable[6][73] ) );
  LHQD1BWP \vrf/regTable_reg[6][74]  ( .E(n5139), .D(\vrf/N92 ), .Q(
        \vrf/regTable[6][74] ) );
  LHQD1BWP \vrf/regTable_reg[6][75]  ( .E(n5139), .D(\vrf/N93 ), .Q(
        \vrf/regTable[6][75] ) );
  LHQD1BWP \vrf/regTable_reg[6][76]  ( .E(n5139), .D(\vrf/N94 ), .Q(
        \vrf/regTable[6][76] ) );
  LHQD1BWP \vrf/regTable_reg[6][77]  ( .E(n5139), .D(\vrf/N95 ), .Q(
        \vrf/regTable[6][77] ) );
  LHQD1BWP \vrf/regTable_reg[6][78]  ( .E(n5139), .D(\vrf/N96 ), .Q(
        \vrf/regTable[6][78] ) );
  LHQD1BWP \vrf/regTable_reg[6][79]  ( .E(n5138), .D(\vrf/N97 ), .Q(
        \vrf/regTable[6][79] ) );
  LHQD1BWP \vrf/regTable_reg[6][80]  ( .E(n5138), .D(\vrf/N98 ), .Q(
        \vrf/regTable[6][80] ) );
  LHQD1BWP \vrf/regTable_reg[6][81]  ( .E(n5138), .D(\vrf/N99 ), .Q(
        \vrf/regTable[6][81] ) );
  LHQD1BWP \vrf/regTable_reg[6][82]  ( .E(n5138), .D(\vrf/N100 ), .Q(
        \vrf/regTable[6][82] ) );
  LHQD1BWP \vrf/regTable_reg[6][83]  ( .E(n5138), .D(\vrf/N101 ), .Q(
        \vrf/regTable[6][83] ) );
  LHQD1BWP \vrf/regTable_reg[6][84]  ( .E(n5138), .D(\vrf/N102 ), .Q(
        \vrf/regTable[6][84] ) );
  LHQD1BWP \vrf/regTable_reg[6][85]  ( .E(n5138), .D(\vrf/N103 ), .Q(
        \vrf/regTable[6][85] ) );
  LHQD1BWP \vrf/regTable_reg[6][86]  ( .E(n5138), .D(\vrf/N104 ), .Q(
        \vrf/regTable[6][86] ) );
  LHQD1BWP \vrf/regTable_reg[6][87]  ( .E(n5138), .D(\vrf/N105 ), .Q(
        \vrf/regTable[6][87] ) );
  LHQD1BWP \vrf/regTable_reg[6][88]  ( .E(n5138), .D(\vrf/N106 ), .Q(
        \vrf/regTable[6][88] ) );
  LHQD1BWP \vrf/regTable_reg[6][89]  ( .E(n5138), .D(\vrf/N107 ), .Q(
        \vrf/regTable[6][89] ) );
  LHQD1BWP \vrf/regTable_reg[6][90]  ( .E(n5137), .D(\vrf/N108 ), .Q(
        \vrf/regTable[6][90] ) );
  LHQD1BWP \vrf/regTable_reg[6][91]  ( .E(n5137), .D(\vrf/N109 ), .Q(
        \vrf/regTable[6][91] ) );
  LHQD1BWP \vrf/regTable_reg[6][92]  ( .E(n5137), .D(\vrf/N110 ), .Q(
        \vrf/regTable[6][92] ) );
  LHQD1BWP \vrf/regTable_reg[6][93]  ( .E(n5137), .D(\vrf/N111 ), .Q(
        \vrf/regTable[6][93] ) );
  LHQD1BWP \vrf/regTable_reg[6][94]  ( .E(n5137), .D(\vrf/N112 ), .Q(
        \vrf/regTable[6][94] ) );
  LHQD1BWP \vrf/regTable_reg[6][95]  ( .E(n5137), .D(\vrf/N113 ), .Q(
        \vrf/regTable[6][95] ) );
  LHQD1BWP \vrf/regTable_reg[6][96]  ( .E(n5137), .D(\vrf/N114 ), .Q(
        \vrf/regTable[6][96] ) );
  LHQD1BWP \vrf/regTable_reg[6][97]  ( .E(n5137), .D(\vrf/N115 ), .Q(
        \vrf/regTable[6][97] ) );
  LHQD1BWP \vrf/regTable_reg[6][98]  ( .E(n5137), .D(\vrf/N116 ), .Q(
        \vrf/regTable[6][98] ) );
  LHQD1BWP \vrf/regTable_reg[6][99]  ( .E(n5137), .D(\vrf/N118 ), .Q(
        \vrf/regTable[6][99] ) );
  LHQD1BWP \vrf/regTable_reg[6][100]  ( .E(n5147), .D(\vrf/N119 ), .Q(
        \vrf/regTable[6][100] ) );
  LHQD1BWP \vrf/regTable_reg[6][101]  ( .E(n5147), .D(\vrf/N120 ), .Q(
        \vrf/regTable[6][101] ) );
  LHQD1BWP \vrf/regTable_reg[6][102]  ( .E(n5147), .D(\vrf/N121 ), .Q(
        \vrf/regTable[6][102] ) );
  LHQD1BWP \vrf/regTable_reg[6][103]  ( .E(n5147), .D(\vrf/N122 ), .Q(
        \vrf/regTable[6][103] ) );
  LHQD1BWP \vrf/regTable_reg[6][104]  ( .E(n5147), .D(\vrf/N123 ), .Q(
        \vrf/regTable[6][104] ) );
  LHQD1BWP \vrf/regTable_reg[6][105]  ( .E(n5146), .D(\vrf/N124 ), .Q(
        \vrf/regTable[6][105] ) );
  LHQD1BWP \vrf/regTable_reg[6][106]  ( .E(n5146), .D(\vrf/N125 ), .Q(
        \vrf/regTable[6][106] ) );
  LHQD1BWP \vrf/regTable_reg[6][107]  ( .E(n5146), .D(\vrf/N126 ), .Q(
        \vrf/regTable[6][107] ) );
  LHQD1BWP \vrf/regTable_reg[6][108]  ( .E(n5146), .D(\vrf/N127 ), .Q(
        \vrf/regTable[6][108] ) );
  LHQD1BWP \vrf/regTable_reg[6][109]  ( .E(n5146), .D(\vrf/N128 ), .Q(
        \vrf/regTable[6][109] ) );
  LHQD1BWP \vrf/regTable_reg[6][110]  ( .E(n5146), .D(\vrf/N129 ), .Q(
        \vrf/regTable[6][110] ) );
  LHQD1BWP \vrf/regTable_reg[6][111]  ( .E(n5146), .D(\vrf/N130 ), .Q(
        \vrf/regTable[6][111] ) );
  LHQD1BWP \vrf/regTable_reg[6][112]  ( .E(n5146), .D(\vrf/N131 ), .Q(
        \vrf/regTable[6][112] ) );
  LHQD1BWP \vrf/regTable_reg[6][113]  ( .E(n5146), .D(\vrf/N132 ), .Q(
        \vrf/regTable[6][113] ) );
  LHQD1BWP \vrf/regTable_reg[6][114]  ( .E(n5146), .D(\vrf/N133 ), .Q(
        \vrf/regTable[6][114] ) );
  LHQD1BWP \vrf/regTable_reg[6][115]  ( .E(n5146), .D(\vrf/N134 ), .Q(
        \vrf/regTable[6][115] ) );
  LHQD1BWP \vrf/regTable_reg[6][116]  ( .E(n5145), .D(\vrf/N135 ), .Q(
        \vrf/regTable[6][116] ) );
  LHQD1BWP \vrf/regTable_reg[6][117]  ( .E(n5145), .D(\vrf/N136 ), .Q(
        \vrf/regTable[6][117] ) );
  LHQD1BWP \vrf/regTable_reg[6][118]  ( .E(n5145), .D(\vrf/N137 ), .Q(
        \vrf/regTable[6][118] ) );
  LHQD1BWP \vrf/regTable_reg[6][119]  ( .E(n5145), .D(\vrf/N138 ), .Q(
        \vrf/regTable[6][119] ) );
  LHQD1BWP \vrf/regTable_reg[6][120]  ( .E(n5145), .D(\vrf/N139 ), .Q(
        \vrf/regTable[6][120] ) );
  LHQD1BWP \vrf/regTable_reg[6][121]  ( .E(n5145), .D(\vrf/N140 ), .Q(
        \vrf/regTable[6][121] ) );
  LHQD1BWP \vrf/regTable_reg[6][122]  ( .E(n5145), .D(\vrf/N141 ), .Q(
        \vrf/regTable[6][122] ) );
  LHQD1BWP \vrf/regTable_reg[6][123]  ( .E(n5145), .D(\vrf/N142 ), .Q(
        \vrf/regTable[6][123] ) );
  LHQD1BWP \vrf/regTable_reg[6][124]  ( .E(n5145), .D(\vrf/N143 ), .Q(
        \vrf/regTable[6][124] ) );
  LHQD1BWP \vrf/regTable_reg[6][125]  ( .E(n5145), .D(\vrf/N144 ), .Q(
        \vrf/regTable[6][125] ) );
  LHQD1BWP \vrf/regTable_reg[6][126]  ( .E(n5145), .D(\vrf/N145 ), .Q(
        \vrf/regTable[6][126] ) );
  LHQD1BWP \vrf/regTable_reg[6][127]  ( .E(n5144), .D(\vrf/N146 ), .Q(
        \vrf/regTable[6][127] ) );
  LHQD1BWP \vrf/regTable_reg[6][128]  ( .E(n5147), .D(\vrf/N147 ), .Q(
        \vrf/regTable[6][128] ) );
  LHQD1BWP \vrf/regTable_reg[6][129]  ( .E(n5147), .D(\vrf/N148 ), .Q(
        \vrf/regTable[6][129] ) );
  LHQD1BWP \vrf/regTable_reg[6][130]  ( .E(n5147), .D(\vrf/N149 ), .Q(
        \vrf/regTable[6][130] ) );
  LHQD1BWP \vrf/regTable_reg[6][131]  ( .E(n5147), .D(\vrf/N150 ), .Q(
        \vrf/regTable[6][131] ) );
  LHQD1BWP \vrf/regTable_reg[6][132]  ( .E(n5147), .D(\vrf/N151 ), .Q(
        \vrf/regTable[6][132] ) );
  LHQD1BWP \vrf/regTable_reg[6][133]  ( .E(n5147), .D(\vrf/N152 ), .Q(
        \vrf/regTable[6][133] ) );
  LHQD1BWP \vrf/regTable_reg[6][134]  ( .E(n5148), .D(\vrf/N153 ), .Q(
        \vrf/regTable[6][134] ) );
  LHQD1BWP \vrf/regTable_reg[6][135]  ( .E(n5148), .D(\vrf/N154 ), .Q(
        \vrf/regTable[6][135] ) );
  LHQD1BWP \vrf/regTable_reg[6][136]  ( .E(n5148), .D(\vrf/N155 ), .Q(
        \vrf/regTable[6][136] ) );
  LHQD1BWP \vrf/regTable_reg[6][137]  ( .E(n5148), .D(\vrf/N156 ), .Q(
        \vrf/regTable[6][137] ) );
  LHQD1BWP \vrf/regTable_reg[6][138]  ( .E(n5148), .D(\vrf/N157 ), .Q(
        \vrf/regTable[6][138] ) );
  LHQD1BWP \vrf/regTable_reg[6][139]  ( .E(n5148), .D(\vrf/N158 ), .Q(
        \vrf/regTable[6][139] ) );
  LHQD1BWP \vrf/regTable_reg[6][140]  ( .E(n5148), .D(\vrf/N159 ), .Q(
        \vrf/regTable[6][140] ) );
  LHQD1BWP \vrf/regTable_reg[6][141]  ( .E(n5148), .D(\vrf/N160 ), .Q(
        \vrf/regTable[6][141] ) );
  LHQD1BWP \vrf/regTable_reg[6][142]  ( .E(n5148), .D(\vrf/N161 ), .Q(
        \vrf/regTable[6][142] ) );
  LHQD1BWP \vrf/regTable_reg[6][143]  ( .E(n5148), .D(\vrf/N162 ), .Q(
        \vrf/regTable[6][143] ) );
  LHQD1BWP \vrf/regTable_reg[6][144]  ( .E(n5148), .D(\vrf/N163 ), .Q(
        \vrf/regTable[6][144] ) );
  LHQD1BWP \vrf/regTable_reg[6][145]  ( .E(n5148), .D(\vrf/N164 ), .Q(
        \vrf/regTable[6][145] ) );
  LHQD1BWP \vrf/regTable_reg[6][146]  ( .E(n5149), .D(\vrf/N165 ), .Q(
        \vrf/regTable[6][146] ) );
  LHQD1BWP \vrf/regTable_reg[6][147]  ( .E(n5149), .D(\vrf/N166 ), .Q(
        \vrf/regTable[6][147] ) );
  LHQD1BWP \vrf/regTable_reg[6][148]  ( .E(n5149), .D(\vrf/N167 ), .Q(
        \vrf/regTable[6][148] ) );
  LHQD1BWP \vrf/regTable_reg[6][149]  ( .E(n5149), .D(\vrf/N168 ), .Q(
        \vrf/regTable[6][149] ) );
  LHQD1BWP \vrf/regTable_reg[6][150]  ( .E(n5149), .D(\vrf/N169 ), .Q(
        \vrf/regTable[6][150] ) );
  LHQD1BWP \vrf/regTable_reg[6][151]  ( .E(n5149), .D(\vrf/N170 ), .Q(
        \vrf/regTable[6][151] ) );
  LHQD1BWP \vrf/regTable_reg[6][152]  ( .E(n5149), .D(\vrf/N171 ), .Q(
        \vrf/regTable[6][152] ) );
  LHQD1BWP \vrf/regTable_reg[6][153]  ( .E(n5149), .D(\vrf/N172 ), .Q(
        \vrf/regTable[6][153] ) );
  LHQD1BWP \vrf/regTable_reg[6][154]  ( .E(n5149), .D(\vrf/N173 ), .Q(
        \vrf/regTable[6][154] ) );
  LHQD1BWP \vrf/regTable_reg[6][155]  ( .E(n5149), .D(\vrf/N174 ), .Q(
        \vrf/regTable[6][155] ) );
  LHQD1BWP \vrf/regTable_reg[6][156]  ( .E(n5149), .D(\vrf/N175 ), .Q(
        \vrf/regTable[6][156] ) );
  LHQD1BWP \vrf/regTable_reg[6][157]  ( .E(n5149), .D(\vrf/N176 ), .Q(
        \vrf/regTable[6][157] ) );
  LHQD1BWP \vrf/regTable_reg[6][158]  ( .E(n5150), .D(\vrf/N177 ), .Q(
        \vrf/regTable[6][158] ) );
  LHQD1BWP \vrf/regTable_reg[6][159]  ( .E(n5150), .D(\vrf/N178 ), .Q(
        \vrf/regTable[6][159] ) );
  LHQD1BWP \vrf/regTable_reg[6][160]  ( .E(n5150), .D(\vrf/N179 ), .Q(
        \vrf/regTable[6][160] ) );
  LHQD1BWP \vrf/regTable_reg[6][161]  ( .E(n5150), .D(\vrf/N180 ), .Q(
        \vrf/regTable[6][161] ) );
  LHQD1BWP \vrf/regTable_reg[6][162]  ( .E(n5150), .D(\vrf/N181 ), .Q(
        \vrf/regTable[6][162] ) );
  LHQD1BWP \vrf/regTable_reg[6][163]  ( .E(n5150), .D(\vrf/N182 ), .Q(
        \vrf/regTable[6][163] ) );
  LHQD1BWP \vrf/regTable_reg[6][164]  ( .E(n5150), .D(\vrf/N183 ), .Q(
        \vrf/regTable[6][164] ) );
  LHQD1BWP \vrf/regTable_reg[6][165]  ( .E(n5150), .D(\vrf/N184 ), .Q(
        \vrf/regTable[6][165] ) );
  LHQD1BWP \vrf/regTable_reg[6][166]  ( .E(n5150), .D(\vrf/N185 ), .Q(
        \vrf/regTable[6][166] ) );
  LHQD1BWP \vrf/regTable_reg[6][167]  ( .E(n5150), .D(\vrf/N186 ), .Q(
        \vrf/regTable[6][167] ) );
  LHQD1BWP \vrf/regTable_reg[6][168]  ( .E(n5150), .D(\vrf/N187 ), .Q(
        \vrf/regTable[6][168] ) );
  LHQD1BWP \vrf/regTable_reg[6][169]  ( .E(n5150), .D(\vrf/N188 ), .Q(
        \vrf/regTable[6][169] ) );
  LHQD1BWP \vrf/regTable_reg[6][170]  ( .E(n5151), .D(\vrf/N189 ), .Q(
        \vrf/regTable[6][170] ) );
  LHQD1BWP \vrf/regTable_reg[6][171]  ( .E(n5151), .D(\vrf/N190 ), .Q(
        \vrf/regTable[6][171] ) );
  LHQD1BWP \vrf/regTable_reg[6][172]  ( .E(n5151), .D(\vrf/N191 ), .Q(
        \vrf/regTable[6][172] ) );
  LHQD1BWP \vrf/regTable_reg[6][173]  ( .E(n5151), .D(\vrf/N192 ), .Q(
        \vrf/regTable[6][173] ) );
  LHQD1BWP \vrf/regTable_reg[6][174]  ( .E(n5151), .D(\vrf/N193 ), .Q(
        \vrf/regTable[6][174] ) );
  LHQD1BWP \vrf/regTable_reg[6][175]  ( .E(n5151), .D(\vrf/N194 ), .Q(
        \vrf/regTable[6][175] ) );
  LHQD1BWP \vrf/regTable_reg[6][176]  ( .E(n5151), .D(\vrf/N195 ), .Q(
        \vrf/regTable[6][176] ) );
  LHQD1BWP \vrf/regTable_reg[6][177]  ( .E(n5151), .D(\vrf/N196 ), .Q(
        \vrf/regTable[6][177] ) );
  LHQD1BWP \vrf/regTable_reg[6][178]  ( .E(n5151), .D(\vrf/N197 ), .Q(
        \vrf/regTable[6][178] ) );
  LHQD1BWP \vrf/regTable_reg[6][179]  ( .E(n5151), .D(\vrf/N198 ), .Q(
        \vrf/regTable[6][179] ) );
  LHQD1BWP \vrf/regTable_reg[6][180]  ( .E(n5151), .D(\vrf/N199 ), .Q(
        \vrf/regTable[6][180] ) );
  LHQD1BWP \vrf/regTable_reg[6][181]  ( .E(n5151), .D(\vrf/N200 ), .Q(
        \vrf/regTable[6][181] ) );
  LHQD1BWP \vrf/regTable_reg[6][182]  ( .E(n5152), .D(\vrf/N201 ), .Q(
        \vrf/regTable[6][182] ) );
  LHQD1BWP \vrf/regTable_reg[6][183]  ( .E(n5152), .D(\vrf/N202 ), .Q(
        \vrf/regTable[6][183] ) );
  LHQD1BWP \vrf/regTable_reg[6][184]  ( .E(n5152), .D(\vrf/N203 ), .Q(
        \vrf/regTable[6][184] ) );
  LHQD1BWP \vrf/regTable_reg[6][185]  ( .E(n5152), .D(\vrf/N204 ), .Q(
        \vrf/regTable[6][185] ) );
  LHQD1BWP \vrf/regTable_reg[6][186]  ( .E(n5152), .D(\vrf/N205 ), .Q(
        \vrf/regTable[6][186] ) );
  LHQD1BWP \vrf/regTable_reg[6][187]  ( .E(n5152), .D(\vrf/N206 ), .Q(
        \vrf/regTable[6][187] ) );
  LHQD1BWP \vrf/regTable_reg[6][188]  ( .E(n5152), .D(\vrf/N207 ), .Q(
        \vrf/regTable[6][188] ) );
  LHQD1BWP \vrf/regTable_reg[6][189]  ( .E(n5152), .D(\vrf/N208 ), .Q(
        \vrf/regTable[6][189] ) );
  LHQD1BWP \vrf/regTable_reg[6][190]  ( .E(n5152), .D(\vrf/N209 ), .Q(
        \vrf/regTable[6][190] ) );
  LHQD1BWP \vrf/regTable_reg[6][191]  ( .E(n5152), .D(\vrf/N210 ), .Q(
        \vrf/regTable[6][191] ) );
  LHQD1BWP \vrf/regTable_reg[6][192]  ( .E(n5152), .D(\vrf/N211 ), .Q(
        \vrf/regTable[6][192] ) );
  LHQD1BWP \vrf/regTable_reg[6][193]  ( .E(n5152), .D(\vrf/N212 ), .Q(
        \vrf/regTable[6][193] ) );
  LHQD1BWP \vrf/regTable_reg[6][194]  ( .E(n5153), .D(\vrf/N213 ), .Q(
        \vrf/regTable[6][194] ) );
  LHQD1BWP \vrf/regTable_reg[6][195]  ( .E(n5153), .D(\vrf/N214 ), .Q(
        \vrf/regTable[6][195] ) );
  LHQD1BWP \vrf/regTable_reg[6][196]  ( .E(n5153), .D(\vrf/N215 ), .Q(
        \vrf/regTable[6][196] ) );
  LHQD1BWP \vrf/regTable_reg[6][197]  ( .E(n5153), .D(\vrf/N216 ), .Q(
        \vrf/regTable[6][197] ) );
  LHQD1BWP \vrf/regTable_reg[6][198]  ( .E(n5153), .D(\vrf/N218 ), .Q(
        \vrf/regTable[6][198] ) );
  LHQD1BWP \vrf/regTable_reg[6][199]  ( .E(n5153), .D(\vrf/N219 ), .Q(
        \vrf/regTable[6][199] ) );
  LHQD1BWP \vrf/regTable_reg[6][200]  ( .E(n5153), .D(\vrf/N220 ), .Q(
        \vrf/regTable[6][200] ) );
  LHQD1BWP \vrf/regTable_reg[6][201]  ( .E(n5153), .D(\vrf/N221 ), .Q(
        \vrf/regTable[6][201] ) );
  LHQD1BWP \vrf/regTable_reg[6][202]  ( .E(n5153), .D(\vrf/N222 ), .Q(
        \vrf/regTable[6][202] ) );
  LHQD1BWP \vrf/regTable_reg[6][203]  ( .E(n5153), .D(\vrf/N223 ), .Q(
        \vrf/regTable[6][203] ) );
  LHQD1BWP \vrf/regTable_reg[6][204]  ( .E(n5153), .D(\vrf/N224 ), .Q(
        \vrf/regTable[6][204] ) );
  LHQD1BWP \vrf/regTable_reg[6][205]  ( .E(n5153), .D(\vrf/N225 ), .Q(
        \vrf/regTable[6][205] ) );
  LHQD1BWP \vrf/regTable_reg[6][206]  ( .E(n5154), .D(\vrf/N226 ), .Q(
        \vrf/regTable[6][206] ) );
  LHQD1BWP \vrf/regTable_reg[6][207]  ( .E(n5154), .D(\vrf/N227 ), .Q(
        \vrf/regTable[6][207] ) );
  LHQD1BWP \vrf/regTable_reg[6][208]  ( .E(n5154), .D(\vrf/N228 ), .Q(
        \vrf/regTable[6][208] ) );
  LHQD1BWP \vrf/regTable_reg[6][209]  ( .E(n5154), .D(\vrf/N229 ), .Q(
        \vrf/regTable[6][209] ) );
  LHQD1BWP \vrf/regTable_reg[6][210]  ( .E(n5154), .D(\vrf/N230 ), .Q(
        \vrf/regTable[6][210] ) );
  LHQD1BWP \vrf/regTable_reg[6][211]  ( .E(n5154), .D(\vrf/N231 ), .Q(
        \vrf/regTable[6][211] ) );
  LHQD1BWP \vrf/regTable_reg[6][212]  ( .E(n5154), .D(\vrf/N232 ), .Q(
        \vrf/regTable[6][212] ) );
  LHQD1BWP \vrf/regTable_reg[6][213]  ( .E(n5154), .D(\vrf/N233 ), .Q(
        \vrf/regTable[6][213] ) );
  LHQD1BWP \vrf/regTable_reg[6][214]  ( .E(n5154), .D(\vrf/N234 ), .Q(
        \vrf/regTable[6][214] ) );
  LHQD1BWP \vrf/regTable_reg[6][215]  ( .E(n5154), .D(\vrf/N235 ), .Q(
        \vrf/regTable[6][215] ) );
  LHQD1BWP \vrf/regTable_reg[6][216]  ( .E(n5154), .D(\vrf/N236 ), .Q(
        \vrf/regTable[6][216] ) );
  LHQD1BWP \vrf/regTable_reg[6][217]  ( .E(n5154), .D(\vrf/N237 ), .Q(
        \vrf/regTable[6][217] ) );
  LHQD1BWP \vrf/regTable_reg[6][218]  ( .E(n5155), .D(\vrf/N238 ), .Q(
        \vrf/regTable[6][218] ) );
  LHQD1BWP \vrf/regTable_reg[6][219]  ( .E(n5155), .D(\vrf/N239 ), .Q(
        \vrf/regTable[6][219] ) );
  LHQD1BWP \vrf/regTable_reg[6][220]  ( .E(n5155), .D(\vrf/N240 ), .Q(
        \vrf/regTable[6][220] ) );
  LHQD1BWP \vrf/regTable_reg[6][221]  ( .E(n5155), .D(\vrf/N241 ), .Q(
        \vrf/regTable[6][221] ) );
  LHQD1BWP \vrf/regTable_reg[6][222]  ( .E(n5155), .D(\vrf/N242 ), .Q(
        \vrf/regTable[6][222] ) );
  LHQD1BWP \vrf/regTable_reg[6][223]  ( .E(n5155), .D(\vrf/N243 ), .Q(
        \vrf/regTable[6][223] ) );
  LHQD1BWP \vrf/regTable_reg[6][224]  ( .E(n5155), .D(\vrf/N244 ), .Q(
        \vrf/regTable[6][224] ) );
  LHQD1BWP \vrf/regTable_reg[6][225]  ( .E(n5155), .D(\vrf/N245 ), .Q(
        \vrf/regTable[6][225] ) );
  LHQD1BWP \vrf/regTable_reg[6][226]  ( .E(n5155), .D(\vrf/N246 ), .Q(
        \vrf/regTable[6][226] ) );
  LHQD1BWP \vrf/regTable_reg[6][227]  ( .E(n5155), .D(\vrf/N247 ), .Q(
        \vrf/regTable[6][227] ) );
  LHQD1BWP \vrf/regTable_reg[6][228]  ( .E(n5155), .D(\vrf/N248 ), .Q(
        \vrf/regTable[6][228] ) );
  LHQD1BWP \vrf/regTable_reg[6][229]  ( .E(n5155), .D(\vrf/N249 ), .Q(
        \vrf/regTable[6][229] ) );
  LHQD1BWP \vrf/regTable_reg[6][230]  ( .E(n5156), .D(\vrf/N250 ), .Q(
        \vrf/regTable[6][230] ) );
  LHQD1BWP \vrf/regTable_reg[6][231]  ( .E(n5156), .D(\vrf/N251 ), .Q(
        \vrf/regTable[6][231] ) );
  LHQD1BWP \vrf/regTable_reg[6][232]  ( .E(n5156), .D(\vrf/N252 ), .Q(
        \vrf/regTable[6][232] ) );
  LHQD1BWP \vrf/regTable_reg[6][233]  ( .E(n5156), .D(\vrf/N253 ), .Q(
        \vrf/regTable[6][233] ) );
  LHQD1BWP \vrf/regTable_reg[6][234]  ( .E(n5156), .D(\vrf/N254 ), .Q(
        \vrf/regTable[6][234] ) );
  LHQD1BWP \vrf/regTable_reg[6][235]  ( .E(n5156), .D(\vrf/N255 ), .Q(
        \vrf/regTable[6][235] ) );
  LHQD1BWP \vrf/regTable_reg[6][236]  ( .E(n5156), .D(\vrf/N256 ), .Q(
        \vrf/regTable[6][236] ) );
  LHQD1BWP \vrf/regTable_reg[6][237]  ( .E(n5156), .D(\vrf/N257 ), .Q(
        \vrf/regTable[6][237] ) );
  LHQD1BWP \vrf/regTable_reg[6][238]  ( .E(n5156), .D(\vrf/N258 ), .Q(
        \vrf/regTable[6][238] ) );
  LHQD1BWP \vrf/regTable_reg[6][239]  ( .E(n5156), .D(\vrf/N259 ), .Q(
        \vrf/regTable[6][239] ) );
  LHQD1BWP \vrf/regTable_reg[6][240]  ( .E(n5156), .D(\vrf/N260 ), .Q(
        \vrf/regTable[6][240] ) );
  LHQD1BWP \vrf/regTable_reg[6][241]  ( .E(n5156), .D(\vrf/N261 ), .Q(
        \vrf/regTable[6][241] ) );
  LHQD1BWP \vrf/regTable_reg[6][242]  ( .E(n5157), .D(\vrf/N262 ), .Q(
        \vrf/regTable[6][242] ) );
  LHQD1BWP \vrf/regTable_reg[6][243]  ( .E(n5157), .D(\vrf/N263 ), .Q(
        \vrf/regTable[6][243] ) );
  LHQD1BWP \vrf/regTable_reg[6][244]  ( .E(n5157), .D(\vrf/N264 ), .Q(
        \vrf/regTable[6][244] ) );
  LHQD1BWP \vrf/regTable_reg[6][245]  ( .E(n5157), .D(\vrf/N265 ), .Q(
        \vrf/regTable[6][245] ) );
  LHQD1BWP \vrf/regTable_reg[6][246]  ( .E(n5157), .D(\vrf/N266 ), .Q(
        \vrf/regTable[6][246] ) );
  LHQD1BWP \vrf/regTable_reg[6][247]  ( .E(n5157), .D(\vrf/N267 ), .Q(
        \vrf/regTable[6][247] ) );
  LHQD1BWP \vrf/regTable_reg[6][248]  ( .E(n5157), .D(\vrf/N268 ), .Q(
        \vrf/regTable[6][248] ) );
  LHQD1BWP \vrf/regTable_reg[6][249]  ( .E(n5157), .D(\vrf/N269 ), .Q(
        \vrf/regTable[6][249] ) );
  LHQD1BWP \vrf/regTable_reg[6][250]  ( .E(n5157), .D(\vrf/N270 ), .Q(
        \vrf/regTable[6][250] ) );
  LHQD1BWP \vrf/regTable_reg[6][251]  ( .E(n5157), .D(\vrf/N271 ), .Q(
        \vrf/regTable[6][251] ) );
  LHQD1BWP \vrf/regTable_reg[6][252]  ( .E(n5157), .D(\vrf/N272 ), .Q(
        \vrf/regTable[6][252] ) );
  LHQD1BWP \vrf/regTable_reg[6][253]  ( .E(n5157), .D(\vrf/N273 ), .Q(
        \vrf/regTable[6][253] ) );
  LHQD1BWP \vrf/regTable_reg[2][0]  ( .E(n5283), .D(\vrf/N18 ), .Q(
        \vrf/regTable[2][0] ) );
  LHQD1BWP \vrf/regTable_reg[2][1]  ( .E(n5280), .D(\vrf/N19 ), .Q(
        \vrf/regTable[2][1] ) );
  LHQD1BWP \vrf/regTable_reg[2][2]  ( .E(n5279), .D(\vrf/N20 ), .Q(
        \vrf/regTable[2][2] ) );
  LHQD1BWP \vrf/regTable_reg[2][3]  ( .E(n5278), .D(\vrf/N21 ), .Q(
        \vrf/regTable[2][3] ) );
  LHQD1BWP \vrf/regTable_reg[2][4]  ( .E(n5277), .D(\vrf/N22 ), .Q(
        \vrf/regTable[2][4] ) );
  LHQD1BWP \vrf/regTable_reg[2][5]  ( .E(n5276), .D(\vrf/N23 ), .Q(
        \vrf/regTable[2][5] ) );
  LHQD1BWP \vrf/regTable_reg[2][6]  ( .E(n5275), .D(\vrf/N24 ), .Q(
        \vrf/regTable[2][6] ) );
  LHQD1BWP \vrf/regTable_reg[2][7]  ( .E(n5274), .D(\vrf/N25 ), .Q(
        \vrf/regTable[2][7] ) );
  LHQD1BWP \vrf/regTable_reg[2][8]  ( .E(n5273), .D(\vrf/N26 ), .Q(
        \vrf/regTable[2][8] ) );
  LHQD1BWP \vrf/regTable_reg[2][9]  ( .E(n5273), .D(\vrf/N27 ), .Q(
        \vrf/regTable[2][9] ) );
  LHQD1BWP \vrf/regTable_reg[2][10]  ( .E(n5282), .D(\vrf/N28 ), .Q(
        \vrf/regTable[2][10] ) );
  LHQD1BWP \vrf/regTable_reg[2][11]  ( .E(n5281), .D(\vrf/N29 ), .Q(
        \vrf/regTable[2][11] ) );
  LHQD1BWP \vrf/regTable_reg[2][12]  ( .E(n5280), .D(\vrf/N30 ), .Q(
        \vrf/regTable[2][12] ) );
  LHQD1BWP \vrf/regTable_reg[2][13]  ( .E(n5280), .D(\vrf/N31 ), .Q(
        \vrf/regTable[2][13] ) );
  LHQD1BWP \vrf/regTable_reg[2][14]  ( .E(n5280), .D(\vrf/N32 ), .Q(
        \vrf/regTable[2][14] ) );
  LHQD1BWP \vrf/regTable_reg[2][17]  ( .E(n5280), .D(\vrf/N35 ), .Q(
        \vrf/regTable[2][17] ) );
  LHQD1BWP \vrf/regTable_reg[2][18]  ( .E(n5280), .D(\vrf/N36 ), .Q(
        \vrf/regTable[2][18] ) );
  LHQD1BWP \vrf/regTable_reg[2][19]  ( .E(n5280), .D(\vrf/N37 ), .Q(
        \vrf/regTable[2][19] ) );
  LHQD1BWP \vrf/regTable_reg[2][20]  ( .E(n5280), .D(\vrf/N38 ), .Q(
        \vrf/regTable[2][20] ) );
  LHQD1BWP \vrf/regTable_reg[2][21]  ( .E(n5280), .D(\vrf/N39 ), .Q(
        \vrf/regTable[2][21] ) );
  LHQD1BWP \vrf/regTable_reg[2][22]  ( .E(n5280), .D(\vrf/N40 ), .Q(
        \vrf/regTable[2][22] ) );
  LHQD1BWP \vrf/regTable_reg[2][23]  ( .E(n5280), .D(\vrf/N41 ), .Q(
        \vrf/regTable[2][23] ) );
  LHQD1BWP \vrf/regTable_reg[2][24]  ( .E(n5279), .D(\vrf/N42 ), .Q(
        \vrf/regTable[2][24] ) );
  LHQD1BWP \vrf/regTable_reg[2][25]  ( .E(n5279), .D(\vrf/N43 ), .Q(
        \vrf/regTable[2][25] ) );
  LHQD1BWP \vrf/regTable_reg[2][26]  ( .E(n5279), .D(\vrf/N44 ), .Q(
        \vrf/regTable[2][26] ) );
  LHQD1BWP \vrf/regTable_reg[2][27]  ( .E(n5279), .D(\vrf/N45 ), .Q(
        \vrf/regTable[2][27] ) );
  LHQD1BWP \vrf/regTable_reg[2][28]  ( .E(n5279), .D(\vrf/N46 ), .Q(
        \vrf/regTable[2][28] ) );
  LHQD1BWP \vrf/regTable_reg[2][29]  ( .E(n5279), .D(\vrf/N47 ), .Q(
        \vrf/regTable[2][29] ) );
  LHQD1BWP \vrf/regTable_reg[2][30]  ( .E(n5279), .D(\vrf/N48 ), .Q(
        \vrf/regTable[2][30] ) );
  LHQD1BWP \vrf/regTable_reg[2][31]  ( .E(n5279), .D(\vrf/N49 ), .Q(
        \vrf/regTable[2][31] ) );
  LHQD1BWP \vrf/regTable_reg[2][32]  ( .E(n5279), .D(\vrf/N50 ), .Q(
        \vrf/regTable[2][32] ) );
  LHQD1BWP \vrf/regTable_reg[2][33]  ( .E(n5279), .D(\vrf/N51 ), .Q(
        \vrf/regTable[2][33] ) );
  LHQD1BWP \vrf/regTable_reg[2][34]  ( .E(n5279), .D(\vrf/N52 ), .Q(
        \vrf/regTable[2][34] ) );
  LHQD1BWP \vrf/regTable_reg[2][35]  ( .E(n5278), .D(\vrf/N53 ), .Q(
        \vrf/regTable[2][35] ) );
  LHQD1BWP \vrf/regTable_reg[2][36]  ( .E(n5278), .D(\vrf/N54 ), .Q(
        \vrf/regTable[2][36] ) );
  LHQD1BWP \vrf/regTable_reg[2][37]  ( .E(n5278), .D(\vrf/N55 ), .Q(
        \vrf/regTable[2][37] ) );
  LHQD1BWP \vrf/regTable_reg[2][38]  ( .E(n5278), .D(\vrf/N56 ), .Q(
        \vrf/regTable[2][38] ) );
  LHQD1BWP \vrf/regTable_reg[2][39]  ( .E(n5278), .D(\vrf/N57 ), .Q(
        \vrf/regTable[2][39] ) );
  LHQD1BWP \vrf/regTable_reg[2][40]  ( .E(n5278), .D(\vrf/N58 ), .Q(
        \vrf/regTable[2][40] ) );
  LHQD1BWP \vrf/regTable_reg[2][41]  ( .E(n5278), .D(\vrf/N59 ), .Q(
        \vrf/regTable[2][41] ) );
  LHQD1BWP \vrf/regTable_reg[2][42]  ( .E(n5278), .D(\vrf/N60 ), .Q(
        \vrf/regTable[2][42] ) );
  LHQD1BWP \vrf/regTable_reg[2][43]  ( .E(n5278), .D(\vrf/N61 ), .Q(
        \vrf/regTable[2][43] ) );
  LHQD1BWP \vrf/regTable_reg[2][44]  ( .E(n5278), .D(\vrf/N62 ), .Q(
        \vrf/regTable[2][44] ) );
  LHQD1BWP \vrf/regTable_reg[2][45]  ( .E(n5278), .D(\vrf/N63 ), .Q(
        \vrf/regTable[2][45] ) );
  LHQD1BWP \vrf/regTable_reg[2][46]  ( .E(n5277), .D(\vrf/N64 ), .Q(
        \vrf/regTable[2][46] ) );
  LHQD1BWP \vrf/regTable_reg[2][47]  ( .E(n5277), .D(\vrf/N65 ), .Q(
        \vrf/regTable[2][47] ) );
  LHQD1BWP \vrf/regTable_reg[2][48]  ( .E(n5277), .D(\vrf/N66 ), .Q(
        \vrf/regTable[2][48] ) );
  LHQD1BWP \vrf/regTable_reg[2][49]  ( .E(n5277), .D(\vrf/N67 ), .Q(
        \vrf/regTable[2][49] ) );
  LHQD1BWP \vrf/regTable_reg[2][50]  ( .E(n5277), .D(\vrf/N68 ), .Q(
        \vrf/regTable[2][50] ) );
  LHQD1BWP \vrf/regTable_reg[2][51]  ( .E(n5277), .D(\vrf/N69 ), .Q(
        \vrf/regTable[2][51] ) );
  LHQD1BWP \vrf/regTable_reg[2][52]  ( .E(n5277), .D(\vrf/N70 ), .Q(
        \vrf/regTable[2][52] ) );
  LHQD1BWP \vrf/regTable_reg[2][53]  ( .E(n5277), .D(\vrf/N71 ), .Q(
        \vrf/regTable[2][53] ) );
  LHQD1BWP \vrf/regTable_reg[2][54]  ( .E(n5277), .D(\vrf/N72 ), .Q(
        \vrf/regTable[2][54] ) );
  LHQD1BWP \vrf/regTable_reg[2][55]  ( .E(n5277), .D(\vrf/N73 ), .Q(
        \vrf/regTable[2][55] ) );
  LHQD1BWP \vrf/regTable_reg[2][56]  ( .E(n5277), .D(\vrf/N74 ), .Q(
        \vrf/regTable[2][56] ) );
  LHQD1BWP \vrf/regTable_reg[2][57]  ( .E(n5276), .D(\vrf/N75 ), .Q(
        \vrf/regTable[2][57] ) );
  LHQD1BWP \vrf/regTable_reg[2][58]  ( .E(n5276), .D(\vrf/N76 ), .Q(
        \vrf/regTable[2][58] ) );
  LHQD1BWP \vrf/regTable_reg[2][59]  ( .E(n5276), .D(\vrf/N77 ), .Q(
        \vrf/regTable[2][59] ) );
  LHQD1BWP \vrf/regTable_reg[2][60]  ( .E(n5276), .D(\vrf/N78 ), .Q(
        \vrf/regTable[2][60] ) );
  LHQD1BWP \vrf/regTable_reg[2][61]  ( .E(n5276), .D(\vrf/N79 ), .Q(
        \vrf/regTable[2][61] ) );
  LHQD1BWP \vrf/regTable_reg[2][62]  ( .E(n5276), .D(\vrf/N80 ), .Q(
        \vrf/regTable[2][62] ) );
  LHQD1BWP \vrf/regTable_reg[2][63]  ( .E(n5276), .D(\vrf/N81 ), .Q(
        \vrf/regTable[2][63] ) );
  LHQD1BWP \vrf/regTable_reg[2][64]  ( .E(n5276), .D(\vrf/N82 ), .Q(
        \vrf/regTable[2][64] ) );
  LHQD1BWP \vrf/regTable_reg[2][65]  ( .E(n5276), .D(\vrf/N83 ), .Q(
        \vrf/regTable[2][65] ) );
  LHQD1BWP \vrf/regTable_reg[2][66]  ( .E(n5276), .D(\vrf/N84 ), .Q(
        \vrf/regTable[2][66] ) );
  LHQD1BWP \vrf/regTable_reg[2][67]  ( .E(n5276), .D(\vrf/N85 ), .Q(
        \vrf/regTable[2][67] ) );
  LHQD1BWP \vrf/regTable_reg[2][68]  ( .E(n5275), .D(\vrf/N86 ), .Q(
        \vrf/regTable[2][68] ) );
  LHQD1BWP \vrf/regTable_reg[2][69]  ( .E(n5275), .D(\vrf/N87 ), .Q(
        \vrf/regTable[2][69] ) );
  LHQD1BWP \vrf/regTable_reg[2][70]  ( .E(n5275), .D(\vrf/N88 ), .Q(
        \vrf/regTable[2][70] ) );
  LHQD1BWP \vrf/regTable_reg[2][71]  ( .E(n5275), .D(\vrf/N89 ), .Q(
        \vrf/regTable[2][71] ) );
  LHQD1BWP \vrf/regTable_reg[2][72]  ( .E(n5275), .D(\vrf/N90 ), .Q(
        \vrf/regTable[2][72] ) );
  LHQD1BWP \vrf/regTable_reg[2][73]  ( .E(n5275), .D(\vrf/N91 ), .Q(
        \vrf/regTable[2][73] ) );
  LHQD1BWP \vrf/regTable_reg[2][74]  ( .E(n5275), .D(\vrf/N92 ), .Q(
        \vrf/regTable[2][74] ) );
  LHQD1BWP \vrf/regTable_reg[2][75]  ( .E(n5275), .D(\vrf/N93 ), .Q(
        \vrf/regTable[2][75] ) );
  LHQD1BWP \vrf/regTable_reg[2][76]  ( .E(n5275), .D(\vrf/N94 ), .Q(
        \vrf/regTable[2][76] ) );
  LHQD1BWP \vrf/regTable_reg[2][77]  ( .E(n5275), .D(\vrf/N95 ), .Q(
        \vrf/regTable[2][77] ) );
  LHQD1BWP \vrf/regTable_reg[2][78]  ( .E(n5275), .D(\vrf/N96 ), .Q(
        \vrf/regTable[2][78] ) );
  LHQD1BWP \vrf/regTable_reg[2][79]  ( .E(n5274), .D(\vrf/N97 ), .Q(
        \vrf/regTable[2][79] ) );
  LHQD1BWP \vrf/regTable_reg[2][80]  ( .E(n5274), .D(\vrf/N98 ), .Q(
        \vrf/regTable[2][80] ) );
  LHQD1BWP \vrf/regTable_reg[2][81]  ( .E(n5274), .D(\vrf/N99 ), .Q(
        \vrf/regTable[2][81] ) );
  LHQD1BWP \vrf/regTable_reg[2][82]  ( .E(n5274), .D(\vrf/N100 ), .Q(
        \vrf/regTable[2][82] ) );
  LHQD1BWP \vrf/regTable_reg[2][83]  ( .E(n5274), .D(\vrf/N101 ), .Q(
        \vrf/regTable[2][83] ) );
  LHQD1BWP \vrf/regTable_reg[2][84]  ( .E(n5274), .D(\vrf/N102 ), .Q(
        \vrf/regTable[2][84] ) );
  LHQD1BWP \vrf/regTable_reg[2][85]  ( .E(n5274), .D(\vrf/N103 ), .Q(
        \vrf/regTable[2][85] ) );
  LHQD1BWP \vrf/regTable_reg[2][86]  ( .E(n5274), .D(\vrf/N104 ), .Q(
        \vrf/regTable[2][86] ) );
  LHQD1BWP \vrf/regTable_reg[2][87]  ( .E(n5274), .D(\vrf/N105 ), .Q(
        \vrf/regTable[2][87] ) );
  LHQD1BWP \vrf/regTable_reg[2][88]  ( .E(n5274), .D(\vrf/N106 ), .Q(
        \vrf/regTable[2][88] ) );
  LHQD1BWP \vrf/regTable_reg[2][89]  ( .E(n5274), .D(\vrf/N107 ), .Q(
        \vrf/regTable[2][89] ) );
  LHQD1BWP \vrf/regTable_reg[2][90]  ( .E(n5273), .D(\vrf/N108 ), .Q(
        \vrf/regTable[2][90] ) );
  LHQD1BWP \vrf/regTable_reg[2][91]  ( .E(n5273), .D(\vrf/N109 ), .Q(
        \vrf/regTable[2][91] ) );
  LHQD1BWP \vrf/regTable_reg[2][92]  ( .E(n5273), .D(\vrf/N110 ), .Q(
        \vrf/regTable[2][92] ) );
  LHQD1BWP \vrf/regTable_reg[2][93]  ( .E(n5273), .D(\vrf/N111 ), .Q(
        \vrf/regTable[2][93] ) );
  LHQD1BWP \vrf/regTable_reg[2][94]  ( .E(n5273), .D(\vrf/N112 ), .Q(
        \vrf/regTable[2][94] ) );
  LHQD1BWP \vrf/regTable_reg[2][95]  ( .E(n5273), .D(\vrf/N113 ), .Q(
        \vrf/regTable[2][95] ) );
  LHQD1BWP \vrf/regTable_reg[2][96]  ( .E(n5273), .D(\vrf/N114 ), .Q(
        \vrf/regTable[2][96] ) );
  LHQD1BWP \vrf/regTable_reg[2][97]  ( .E(n5273), .D(\vrf/N115 ), .Q(
        \vrf/regTable[2][97] ) );
  LHQD1BWP \vrf/regTable_reg[2][98]  ( .E(n5273), .D(\vrf/N116 ), .Q(
        \vrf/regTable[2][98] ) );
  LHQD1BWP \vrf/regTable_reg[2][99]  ( .E(n5273), .D(\vrf/N118 ), .Q(
        \vrf/regTable[2][99] ) );
  LHQD1BWP \vrf/regTable_reg[2][100]  ( .E(n5283), .D(\vrf/N119 ), .Q(
        \vrf/regTable[2][100] ) );
  LHQD1BWP \vrf/regTable_reg[2][101]  ( .E(n5283), .D(\vrf/N120 ), .Q(
        \vrf/regTable[2][101] ) );
  LHQD1BWP \vrf/regTable_reg[2][102]  ( .E(n5283), .D(\vrf/N121 ), .Q(
        \vrf/regTable[2][102] ) );
  LHQD1BWP \vrf/regTable_reg[2][103]  ( .E(n5283), .D(\vrf/N122 ), .Q(
        \vrf/regTable[2][103] ) );
  LHQD1BWP \vrf/regTable_reg[2][104]  ( .E(n5283), .D(\vrf/N123 ), .Q(
        \vrf/regTable[2][104] ) );
  LHQD1BWP \vrf/regTable_reg[2][105]  ( .E(n5282), .D(\vrf/N124 ), .Q(
        \vrf/regTable[2][105] ) );
  LHQD1BWP \vrf/regTable_reg[2][106]  ( .E(n5282), .D(\vrf/N125 ), .Q(
        \vrf/regTable[2][106] ) );
  LHQD1BWP \vrf/regTable_reg[2][107]  ( .E(n5282), .D(\vrf/N126 ), .Q(
        \vrf/regTable[2][107] ) );
  LHQD1BWP \vrf/regTable_reg[2][108]  ( .E(n5282), .D(\vrf/N127 ), .Q(
        \vrf/regTable[2][108] ) );
  LHQD1BWP \vrf/regTable_reg[2][109]  ( .E(n5282), .D(\vrf/N128 ), .Q(
        \vrf/regTable[2][109] ) );
  LHQD1BWP \vrf/regTable_reg[2][110]  ( .E(n5282), .D(\vrf/N129 ), .Q(
        \vrf/regTable[2][110] ) );
  LHQD1BWP \vrf/regTable_reg[2][111]  ( .E(n5282), .D(\vrf/N130 ), .Q(
        \vrf/regTable[2][111] ) );
  LHQD1BWP \vrf/regTable_reg[2][112]  ( .E(n5282), .D(\vrf/N131 ), .Q(
        \vrf/regTable[2][112] ) );
  LHQD1BWP \vrf/regTable_reg[2][113]  ( .E(n5282), .D(\vrf/N132 ), .Q(
        \vrf/regTable[2][113] ) );
  LHQD1BWP \vrf/regTable_reg[2][114]  ( .E(n5282), .D(\vrf/N133 ), .Q(
        \vrf/regTable[2][114] ) );
  LHQD1BWP \vrf/regTable_reg[2][115]  ( .E(n5282), .D(\vrf/N134 ), .Q(
        \vrf/regTable[2][115] ) );
  LHQD1BWP \vrf/regTable_reg[2][116]  ( .E(n5281), .D(\vrf/N135 ), .Q(
        \vrf/regTable[2][116] ) );
  LHQD1BWP \vrf/regTable_reg[2][117]  ( .E(n5281), .D(\vrf/N136 ), .Q(
        \vrf/regTable[2][117] ) );
  LHQD1BWP \vrf/regTable_reg[2][118]  ( .E(n5281), .D(\vrf/N137 ), .Q(
        \vrf/regTable[2][118] ) );
  LHQD1BWP \vrf/regTable_reg[2][119]  ( .E(n5281), .D(\vrf/N138 ), .Q(
        \vrf/regTable[2][119] ) );
  LHQD1BWP \vrf/regTable_reg[2][120]  ( .E(n5281), .D(\vrf/N139 ), .Q(
        \vrf/regTable[2][120] ) );
  LHQD1BWP \vrf/regTable_reg[2][121]  ( .E(n5281), .D(\vrf/N140 ), .Q(
        \vrf/regTable[2][121] ) );
  LHQD1BWP \vrf/regTable_reg[2][122]  ( .E(n5281), .D(\vrf/N141 ), .Q(
        \vrf/regTable[2][122] ) );
  LHQD1BWP \vrf/regTable_reg[2][123]  ( .E(n5281), .D(\vrf/N142 ), .Q(
        \vrf/regTable[2][123] ) );
  LHQD1BWP \vrf/regTable_reg[2][124]  ( .E(n5281), .D(\vrf/N143 ), .Q(
        \vrf/regTable[2][124] ) );
  LHQD1BWP \vrf/regTable_reg[2][125]  ( .E(n5281), .D(\vrf/N144 ), .Q(
        \vrf/regTable[2][125] ) );
  LHQD1BWP \vrf/regTable_reg[2][126]  ( .E(n5281), .D(\vrf/N145 ), .Q(
        \vrf/regTable[2][126] ) );
  LHQD1BWP \vrf/regTable_reg[2][127]  ( .E(n5280), .D(\vrf/N146 ), .Q(
        \vrf/regTable[2][127] ) );
  LHQD1BWP \vrf/regTable_reg[2][128]  ( .E(n5283), .D(\vrf/N147 ), .Q(
        \vrf/regTable[2][128] ) );
  LHQD1BWP \vrf/regTable_reg[2][129]  ( .E(n5283), .D(\vrf/N148 ), .Q(
        \vrf/regTable[2][129] ) );
  LHQD1BWP \vrf/regTable_reg[2][130]  ( .E(n5283), .D(\vrf/N149 ), .Q(
        \vrf/regTable[2][130] ) );
  LHQD1BWP \vrf/regTable_reg[2][131]  ( .E(n5283), .D(\vrf/N150 ), .Q(
        \vrf/regTable[2][131] ) );
  LHQD1BWP \vrf/regTable_reg[2][132]  ( .E(n5283), .D(\vrf/N151 ), .Q(
        \vrf/regTable[2][132] ) );
  LHQD1BWP \vrf/regTable_reg[2][133]  ( .E(n5283), .D(\vrf/N152 ), .Q(
        \vrf/regTable[2][133] ) );
  LHQD1BWP \vrf/regTable_reg[2][134]  ( .E(n5284), .D(\vrf/N153 ), .Q(
        \vrf/regTable[2][134] ) );
  LHQD1BWP \vrf/regTable_reg[2][135]  ( .E(n5284), .D(\vrf/N154 ), .Q(
        \vrf/regTable[2][135] ) );
  LHQD1BWP \vrf/regTable_reg[2][136]  ( .E(n5284), .D(\vrf/N155 ), .Q(
        \vrf/regTable[2][136] ) );
  LHQD1BWP \vrf/regTable_reg[2][137]  ( .E(n5284), .D(\vrf/N156 ), .Q(
        \vrf/regTable[2][137] ) );
  LHQD1BWP \vrf/regTable_reg[2][138]  ( .E(n5284), .D(\vrf/N157 ), .Q(
        \vrf/regTable[2][138] ) );
  LHQD1BWP \vrf/regTable_reg[2][139]  ( .E(n5284), .D(\vrf/N158 ), .Q(
        \vrf/regTable[2][139] ) );
  LHQD1BWP \vrf/regTable_reg[2][140]  ( .E(n5284), .D(\vrf/N159 ), .Q(
        \vrf/regTable[2][140] ) );
  LHQD1BWP \vrf/regTable_reg[2][141]  ( .E(n5284), .D(\vrf/N160 ), .Q(
        \vrf/regTable[2][141] ) );
  LHQD1BWP \vrf/regTable_reg[2][142]  ( .E(n5284), .D(\vrf/N161 ), .Q(
        \vrf/regTable[2][142] ) );
  LHQD1BWP \vrf/regTable_reg[2][143]  ( .E(n5284), .D(\vrf/N162 ), .Q(
        \vrf/regTable[2][143] ) );
  LHQD1BWP \vrf/regTable_reg[2][144]  ( .E(n5284), .D(\vrf/N163 ), .Q(
        \vrf/regTable[2][144] ) );
  LHQD1BWP \vrf/regTable_reg[2][145]  ( .E(n5284), .D(\vrf/N164 ), .Q(
        \vrf/regTable[2][145] ) );
  LHQD1BWP \vrf/regTable_reg[2][146]  ( .E(n5285), .D(\vrf/N165 ), .Q(
        \vrf/regTable[2][146] ) );
  LHQD1BWP \vrf/regTable_reg[2][147]  ( .E(n5285), .D(\vrf/N166 ), .Q(
        \vrf/regTable[2][147] ) );
  LHQD1BWP \vrf/regTable_reg[2][148]  ( .E(n5285), .D(\vrf/N167 ), .Q(
        \vrf/regTable[2][148] ) );
  LHQD1BWP \vrf/regTable_reg[2][149]  ( .E(n5285), .D(\vrf/N168 ), .Q(
        \vrf/regTable[2][149] ) );
  LHQD1BWP \vrf/regTable_reg[2][150]  ( .E(n5285), .D(\vrf/N169 ), .Q(
        \vrf/regTable[2][150] ) );
  LHQD1BWP \vrf/regTable_reg[2][151]  ( .E(n5285), .D(\vrf/N170 ), .Q(
        \vrf/regTable[2][151] ) );
  LHQD1BWP \vrf/regTable_reg[2][152]  ( .E(n5285), .D(\vrf/N171 ), .Q(
        \vrf/regTable[2][152] ) );
  LHQD1BWP \vrf/regTable_reg[2][153]  ( .E(n5285), .D(\vrf/N172 ), .Q(
        \vrf/regTable[2][153] ) );
  LHQD1BWP \vrf/regTable_reg[2][154]  ( .E(n5285), .D(\vrf/N173 ), .Q(
        \vrf/regTable[2][154] ) );
  LHQD1BWP \vrf/regTable_reg[2][155]  ( .E(n5285), .D(\vrf/N174 ), .Q(
        \vrf/regTable[2][155] ) );
  LHQD1BWP \vrf/regTable_reg[2][156]  ( .E(n5285), .D(\vrf/N175 ), .Q(
        \vrf/regTable[2][156] ) );
  LHQD1BWP \vrf/regTable_reg[2][157]  ( .E(n5285), .D(\vrf/N176 ), .Q(
        \vrf/regTable[2][157] ) );
  LHQD1BWP \vrf/regTable_reg[2][158]  ( .E(n5286), .D(\vrf/N177 ), .Q(
        \vrf/regTable[2][158] ) );
  LHQD1BWP \vrf/regTable_reg[2][159]  ( .E(n5286), .D(\vrf/N178 ), .Q(
        \vrf/regTable[2][159] ) );
  LHQD1BWP \vrf/regTable_reg[2][160]  ( .E(n5286), .D(\vrf/N179 ), .Q(
        \vrf/regTable[2][160] ) );
  LHQD1BWP \vrf/regTable_reg[2][161]  ( .E(n5286), .D(\vrf/N180 ), .Q(
        \vrf/regTable[2][161] ) );
  LHQD1BWP \vrf/regTable_reg[2][162]  ( .E(n5286), .D(\vrf/N181 ), .Q(
        \vrf/regTable[2][162] ) );
  LHQD1BWP \vrf/regTable_reg[2][163]  ( .E(n5286), .D(\vrf/N182 ), .Q(
        \vrf/regTable[2][163] ) );
  LHQD1BWP \vrf/regTable_reg[2][164]  ( .E(n5286), .D(\vrf/N183 ), .Q(
        \vrf/regTable[2][164] ) );
  LHQD1BWP \vrf/regTable_reg[2][165]  ( .E(n5286), .D(\vrf/N184 ), .Q(
        \vrf/regTable[2][165] ) );
  LHQD1BWP \vrf/regTable_reg[2][166]  ( .E(n5286), .D(\vrf/N185 ), .Q(
        \vrf/regTable[2][166] ) );
  LHQD1BWP \vrf/regTable_reg[2][167]  ( .E(n5286), .D(\vrf/N186 ), .Q(
        \vrf/regTable[2][167] ) );
  LHQD1BWP \vrf/regTable_reg[2][168]  ( .E(n5286), .D(\vrf/N187 ), .Q(
        \vrf/regTable[2][168] ) );
  LHQD1BWP \vrf/regTable_reg[2][169]  ( .E(n5286), .D(\vrf/N188 ), .Q(
        \vrf/regTable[2][169] ) );
  LHQD1BWP \vrf/regTable_reg[2][170]  ( .E(n5287), .D(\vrf/N189 ), .Q(
        \vrf/regTable[2][170] ) );
  LHQD1BWP \vrf/regTable_reg[2][171]  ( .E(n5287), .D(\vrf/N190 ), .Q(
        \vrf/regTable[2][171] ) );
  LHQD1BWP \vrf/regTable_reg[2][172]  ( .E(n5287), .D(\vrf/N191 ), .Q(
        \vrf/regTable[2][172] ) );
  LHQD1BWP \vrf/regTable_reg[2][173]  ( .E(n5287), .D(\vrf/N192 ), .Q(
        \vrf/regTable[2][173] ) );
  LHQD1BWP \vrf/regTable_reg[2][174]  ( .E(n5287), .D(\vrf/N193 ), .Q(
        \vrf/regTable[2][174] ) );
  LHQD1BWP \vrf/regTable_reg[2][175]  ( .E(n5287), .D(\vrf/N194 ), .Q(
        \vrf/regTable[2][175] ) );
  LHQD1BWP \vrf/regTable_reg[2][176]  ( .E(n5287), .D(\vrf/N195 ), .Q(
        \vrf/regTable[2][176] ) );
  LHQD1BWP \vrf/regTable_reg[2][177]  ( .E(n5287), .D(\vrf/N196 ), .Q(
        \vrf/regTable[2][177] ) );
  LHQD1BWP \vrf/regTable_reg[2][178]  ( .E(n5287), .D(\vrf/N197 ), .Q(
        \vrf/regTable[2][178] ) );
  LHQD1BWP \vrf/regTable_reg[2][179]  ( .E(n5287), .D(\vrf/N198 ), .Q(
        \vrf/regTable[2][179] ) );
  LHQD1BWP \vrf/regTable_reg[2][180]  ( .E(n5287), .D(\vrf/N199 ), .Q(
        \vrf/regTable[2][180] ) );
  LHQD1BWP \vrf/regTable_reg[2][181]  ( .E(n5287), .D(\vrf/N200 ), .Q(
        \vrf/regTable[2][181] ) );
  LHQD1BWP \vrf/regTable_reg[2][182]  ( .E(n5288), .D(\vrf/N201 ), .Q(
        \vrf/regTable[2][182] ) );
  LHQD1BWP \vrf/regTable_reg[2][183]  ( .E(n5288), .D(\vrf/N202 ), .Q(
        \vrf/regTable[2][183] ) );
  LHQD1BWP \vrf/regTable_reg[2][184]  ( .E(n5288), .D(\vrf/N203 ), .Q(
        \vrf/regTable[2][184] ) );
  LHQD1BWP \vrf/regTable_reg[2][185]  ( .E(n5288), .D(\vrf/N204 ), .Q(
        \vrf/regTable[2][185] ) );
  LHQD1BWP \vrf/regTable_reg[2][186]  ( .E(n5288), .D(\vrf/N205 ), .Q(
        \vrf/regTable[2][186] ) );
  LHQD1BWP \vrf/regTable_reg[2][187]  ( .E(n5288), .D(\vrf/N206 ), .Q(
        \vrf/regTable[2][187] ) );
  LHQD1BWP \vrf/regTable_reg[2][188]  ( .E(n5288), .D(\vrf/N207 ), .Q(
        \vrf/regTable[2][188] ) );
  LHQD1BWP \vrf/regTable_reg[2][189]  ( .E(n5288), .D(\vrf/N208 ), .Q(
        \vrf/regTable[2][189] ) );
  LHQD1BWP \vrf/regTable_reg[2][190]  ( .E(n5288), .D(\vrf/N209 ), .Q(
        \vrf/regTable[2][190] ) );
  LHQD1BWP \vrf/regTable_reg[2][191]  ( .E(n5288), .D(\vrf/N210 ), .Q(
        \vrf/regTable[2][191] ) );
  LHQD1BWP \vrf/regTable_reg[2][192]  ( .E(n5288), .D(\vrf/N211 ), .Q(
        \vrf/regTable[2][192] ) );
  LHQD1BWP \vrf/regTable_reg[2][193]  ( .E(n5288), .D(\vrf/N212 ), .Q(
        \vrf/regTable[2][193] ) );
  LHQD1BWP \vrf/regTable_reg[2][194]  ( .E(n5289), .D(\vrf/N213 ), .Q(
        \vrf/regTable[2][194] ) );
  LHQD1BWP \vrf/regTable_reg[2][195]  ( .E(n5289), .D(\vrf/N214 ), .Q(
        \vrf/regTable[2][195] ) );
  LHQD1BWP \vrf/regTable_reg[2][196]  ( .E(n5289), .D(\vrf/N215 ), .Q(
        \vrf/regTable[2][196] ) );
  LHQD1BWP \vrf/regTable_reg[2][197]  ( .E(n5289), .D(\vrf/N216 ), .Q(
        \vrf/regTable[2][197] ) );
  LHQD1BWP \vrf/regTable_reg[2][198]  ( .E(n5289), .D(\vrf/N218 ), .Q(
        \vrf/regTable[2][198] ) );
  LHQD1BWP \vrf/regTable_reg[2][199]  ( .E(n5289), .D(\vrf/N219 ), .Q(
        \vrf/regTable[2][199] ) );
  LHQD1BWP \vrf/regTable_reg[2][200]  ( .E(n5289), .D(\vrf/N220 ), .Q(
        \vrf/regTable[2][200] ) );
  LHQD1BWP \vrf/regTable_reg[2][201]  ( .E(n5289), .D(\vrf/N221 ), .Q(
        \vrf/regTable[2][201] ) );
  LHQD1BWP \vrf/regTable_reg[2][202]  ( .E(n5289), .D(\vrf/N222 ), .Q(
        \vrf/regTable[2][202] ) );
  LHQD1BWP \vrf/regTable_reg[2][203]  ( .E(n5289), .D(\vrf/N223 ), .Q(
        \vrf/regTable[2][203] ) );
  LHQD1BWP \vrf/regTable_reg[2][204]  ( .E(n5289), .D(\vrf/N224 ), .Q(
        \vrf/regTable[2][204] ) );
  LHQD1BWP \vrf/regTable_reg[2][205]  ( .E(n5289), .D(\vrf/N225 ), .Q(
        \vrf/regTable[2][205] ) );
  LHQD1BWP \vrf/regTable_reg[2][206]  ( .E(n5290), .D(\vrf/N226 ), .Q(
        \vrf/regTable[2][206] ) );
  LHQD1BWP \vrf/regTable_reg[2][207]  ( .E(n5290), .D(\vrf/N227 ), .Q(
        \vrf/regTable[2][207] ) );
  LHQD1BWP \vrf/regTable_reg[2][208]  ( .E(n5290), .D(\vrf/N228 ), .Q(
        \vrf/regTable[2][208] ) );
  LHQD1BWP \vrf/regTable_reg[2][209]  ( .E(n5290), .D(\vrf/N229 ), .Q(
        \vrf/regTable[2][209] ) );
  LHQD1BWP \vrf/regTable_reg[2][210]  ( .E(n5290), .D(\vrf/N230 ), .Q(
        \vrf/regTable[2][210] ) );
  LHQD1BWP \vrf/regTable_reg[2][211]  ( .E(n5290), .D(\vrf/N231 ), .Q(
        \vrf/regTable[2][211] ) );
  LHQD1BWP \vrf/regTable_reg[2][212]  ( .E(n5290), .D(\vrf/N232 ), .Q(
        \vrf/regTable[2][212] ) );
  LHQD1BWP \vrf/regTable_reg[2][213]  ( .E(n5290), .D(\vrf/N233 ), .Q(
        \vrf/regTable[2][213] ) );
  LHQD1BWP \vrf/regTable_reg[2][214]  ( .E(n5290), .D(\vrf/N234 ), .Q(
        \vrf/regTable[2][214] ) );
  LHQD1BWP \vrf/regTable_reg[2][215]  ( .E(n5290), .D(\vrf/N235 ), .Q(
        \vrf/regTable[2][215] ) );
  LHQD1BWP \vrf/regTable_reg[2][216]  ( .E(n5290), .D(\vrf/N236 ), .Q(
        \vrf/regTable[2][216] ) );
  LHQD1BWP \vrf/regTable_reg[2][217]  ( .E(n5290), .D(\vrf/N237 ), .Q(
        \vrf/regTable[2][217] ) );
  LHQD1BWP \vrf/regTable_reg[2][218]  ( .E(n5291), .D(\vrf/N238 ), .Q(
        \vrf/regTable[2][218] ) );
  LHQD1BWP \vrf/regTable_reg[2][219]  ( .E(n5291), .D(\vrf/N239 ), .Q(
        \vrf/regTable[2][219] ) );
  LHQD1BWP \vrf/regTable_reg[2][220]  ( .E(n5291), .D(\vrf/N240 ), .Q(
        \vrf/regTable[2][220] ) );
  LHQD1BWP \vrf/regTable_reg[2][221]  ( .E(n5291), .D(\vrf/N241 ), .Q(
        \vrf/regTable[2][221] ) );
  LHQD1BWP \vrf/regTable_reg[2][222]  ( .E(n5291), .D(\vrf/N242 ), .Q(
        \vrf/regTable[2][222] ) );
  LHQD1BWP \vrf/regTable_reg[2][223]  ( .E(n5291), .D(\vrf/N243 ), .Q(
        \vrf/regTable[2][223] ) );
  LHQD1BWP \vrf/regTable_reg[2][224]  ( .E(n5291), .D(\vrf/N244 ), .Q(
        \vrf/regTable[2][224] ) );
  LHQD1BWP \vrf/regTable_reg[2][225]  ( .E(n5291), .D(\vrf/N245 ), .Q(
        \vrf/regTable[2][225] ) );
  LHQD1BWP \vrf/regTable_reg[2][226]  ( .E(n5291), .D(\vrf/N246 ), .Q(
        \vrf/regTable[2][226] ) );
  LHQD1BWP \vrf/regTable_reg[2][227]  ( .E(n5291), .D(\vrf/N247 ), .Q(
        \vrf/regTable[2][227] ) );
  LHQD1BWP \vrf/regTable_reg[2][228]  ( .E(n5291), .D(\vrf/N248 ), .Q(
        \vrf/regTable[2][228] ) );
  LHQD1BWP \vrf/regTable_reg[2][229]  ( .E(n5291), .D(\vrf/N249 ), .Q(
        \vrf/regTable[2][229] ) );
  LHQD1BWP \vrf/regTable_reg[2][230]  ( .E(n5292), .D(\vrf/N250 ), .Q(
        \vrf/regTable[2][230] ) );
  LHQD1BWP \vrf/regTable_reg[2][231]  ( .E(n5292), .D(\vrf/N251 ), .Q(
        \vrf/regTable[2][231] ) );
  LHQD1BWP \vrf/regTable_reg[2][232]  ( .E(n5292), .D(\vrf/N252 ), .Q(
        \vrf/regTable[2][232] ) );
  LHQD1BWP \vrf/regTable_reg[2][233]  ( .E(n5292), .D(\vrf/N253 ), .Q(
        \vrf/regTable[2][233] ) );
  LHQD1BWP \vrf/regTable_reg[2][234]  ( .E(n5292), .D(\vrf/N254 ), .Q(
        \vrf/regTable[2][234] ) );
  LHQD1BWP \vrf/regTable_reg[2][235]  ( .E(n5292), .D(\vrf/N255 ), .Q(
        \vrf/regTable[2][235] ) );
  LHQD1BWP \vrf/regTable_reg[2][236]  ( .E(n5292), .D(\vrf/N256 ), .Q(
        \vrf/regTable[2][236] ) );
  LHQD1BWP \vrf/regTable_reg[2][237]  ( .E(n5292), .D(\vrf/N257 ), .Q(
        \vrf/regTable[2][237] ) );
  LHQD1BWP \vrf/regTable_reg[2][238]  ( .E(n5292), .D(\vrf/N258 ), .Q(
        \vrf/regTable[2][238] ) );
  LHQD1BWP \vrf/regTable_reg[2][239]  ( .E(n5292), .D(\vrf/N259 ), .Q(
        \vrf/regTable[2][239] ) );
  LHQD1BWP \vrf/regTable_reg[2][240]  ( .E(n5292), .D(\vrf/N260 ), .Q(
        \vrf/regTable[2][240] ) );
  LHQD1BWP \vrf/regTable_reg[2][241]  ( .E(n5292), .D(\vrf/N261 ), .Q(
        \vrf/regTable[2][241] ) );
  LHQD1BWP \vrf/regTable_reg[2][242]  ( .E(n5293), .D(\vrf/N262 ), .Q(
        \vrf/regTable[2][242] ) );
  LHQD1BWP \vrf/regTable_reg[2][243]  ( .E(n5293), .D(\vrf/N263 ), .Q(
        \vrf/regTable[2][243] ) );
  LHQD1BWP \vrf/regTable_reg[2][244]  ( .E(n5293), .D(\vrf/N264 ), .Q(
        \vrf/regTable[2][244] ) );
  LHQD1BWP \vrf/regTable_reg[2][245]  ( .E(n5293), .D(\vrf/N265 ), .Q(
        \vrf/regTable[2][245] ) );
  LHQD1BWP \vrf/regTable_reg[2][246]  ( .E(n5293), .D(\vrf/N266 ), .Q(
        \vrf/regTable[2][246] ) );
  LHQD1BWP \vrf/regTable_reg[2][247]  ( .E(n5293), .D(\vrf/N267 ), .Q(
        \vrf/regTable[2][247] ) );
  LHQD1BWP \vrf/regTable_reg[2][248]  ( .E(n5293), .D(\vrf/N268 ), .Q(
        \vrf/regTable[2][248] ) );
  LHQD1BWP \vrf/regTable_reg[2][249]  ( .E(n5293), .D(\vrf/N269 ), .Q(
        \vrf/regTable[2][249] ) );
  LHQD1BWP \vrf/regTable_reg[2][250]  ( .E(n5293), .D(\vrf/N270 ), .Q(
        \vrf/regTable[2][250] ) );
  LHQD1BWP \vrf/regTable_reg[2][251]  ( .E(n5293), .D(\vrf/N271 ), .Q(
        \vrf/regTable[2][251] ) );
  LHQD1BWP \vrf/regTable_reg[2][252]  ( .E(n5293), .D(\vrf/N272 ), .Q(
        \vrf/regTable[2][252] ) );
  LHQD1BWP \vrf/regTable_reg[2][253]  ( .E(n5293), .D(\vrf/N273 ), .Q(
        \vrf/regTable[2][253] ) );
  LHQD1BWP \vrf/regTable_reg[4][15]  ( .E(n5226), .D(\vrf/N33 ), .Q(
        \vrf/regTable[4][15] ) );
  LHQD1BWP \vrf/regTable_reg[4][16]  ( .E(n5226), .D(\vrf/N34 ), .Q(
        \vrf/regTable[4][16] ) );
  LHQD1BWP \vrf/regTable_reg[4][254]  ( .E(n5226), .D(\vrf/N274 ), .Q(
        \vrf/regTable[4][254] ) );
  LHQD1BWP \vrf/regTable_reg[4][255]  ( .E(n5226), .D(\vrf/N275 ), .Q(
        \vrf/regTable[4][255] ) );
  LHQD1BWP \vrf/regTable_reg[0][15]  ( .E(n5362), .D(\vrf/N33 ), .Q(
        \vrf/regTable[0][15] ) );
  LHQD1BWP \vrf/regTable_reg[0][16]  ( .E(n5362), .D(\vrf/N34 ), .Q(
        \vrf/regTable[0][16] ) );
  LHQD1BWP \vrf/regTable_reg[0][254]  ( .E(n5362), .D(\vrf/N274 ), .Q(
        \vrf/regTable[0][254] ) );
  LHQD1BWP \vrf/regTable_reg[0][255]  ( .E(n5362), .D(\vrf/N275 ), .Q(
        \vrf/regTable[0][255] ) );
  LHQD1BWP \vrf/regTable_reg[4][0]  ( .E(n5215), .D(\vrf/N18 ), .Q(
        \vrf/regTable[4][0] ) );
  LHQD1BWP \vrf/regTable_reg[4][1]  ( .E(n5212), .D(\vrf/N19 ), .Q(
        \vrf/regTable[4][1] ) );
  LHQD1BWP \vrf/regTable_reg[4][2]  ( .E(n5211), .D(\vrf/N20 ), .Q(
        \vrf/regTable[4][2] ) );
  LHQD1BWP \vrf/regTable_reg[4][3]  ( .E(n5210), .D(\vrf/N21 ), .Q(
        \vrf/regTable[4][3] ) );
  LHQD1BWP \vrf/regTable_reg[4][4]  ( .E(n5209), .D(\vrf/N22 ), .Q(
        \vrf/regTable[4][4] ) );
  LHQD1BWP \vrf/regTable_reg[4][5]  ( .E(n5208), .D(\vrf/N23 ), .Q(
        \vrf/regTable[4][5] ) );
  LHQD1BWP \vrf/regTable_reg[4][6]  ( .E(n5207), .D(\vrf/N24 ), .Q(
        \vrf/regTable[4][6] ) );
  LHQD1BWP \vrf/regTable_reg[4][7]  ( .E(n5206), .D(\vrf/N25 ), .Q(
        \vrf/regTable[4][7] ) );
  LHQD1BWP \vrf/regTable_reg[4][8]  ( .E(n5205), .D(\vrf/N26 ), .Q(
        \vrf/regTable[4][8] ) );
  LHQD1BWP \vrf/regTable_reg[4][9]  ( .E(n5205), .D(\vrf/N27 ), .Q(
        \vrf/regTable[4][9] ) );
  LHQD1BWP \vrf/regTable_reg[4][10]  ( .E(n5214), .D(\vrf/N28 ), .Q(
        \vrf/regTable[4][10] ) );
  LHQD1BWP \vrf/regTable_reg[4][11]  ( .E(n5213), .D(\vrf/N29 ), .Q(
        \vrf/regTable[4][11] ) );
  LHQD1BWP \vrf/regTable_reg[4][12]  ( .E(n5212), .D(\vrf/N30 ), .Q(
        \vrf/regTable[4][12] ) );
  LHQD1BWP \vrf/regTable_reg[4][13]  ( .E(n5212), .D(\vrf/N31 ), .Q(
        \vrf/regTable[4][13] ) );
  LHQD1BWP \vrf/regTable_reg[4][14]  ( .E(n5212), .D(\vrf/N32 ), .Q(
        \vrf/regTable[4][14] ) );
  LHQD1BWP \vrf/regTable_reg[4][17]  ( .E(n5212), .D(\vrf/N35 ), .Q(
        \vrf/regTable[4][17] ) );
  LHQD1BWP \vrf/regTable_reg[4][18]  ( .E(n5212), .D(\vrf/N36 ), .Q(
        \vrf/regTable[4][18] ) );
  LHQD1BWP \vrf/regTable_reg[4][19]  ( .E(n5212), .D(\vrf/N37 ), .Q(
        \vrf/regTable[4][19] ) );
  LHQD1BWP \vrf/regTable_reg[4][20]  ( .E(n5212), .D(\vrf/N38 ), .Q(
        \vrf/regTable[4][20] ) );
  LHQD1BWP \vrf/regTable_reg[4][21]  ( .E(n5212), .D(\vrf/N39 ), .Q(
        \vrf/regTable[4][21] ) );
  LHQD1BWP \vrf/regTable_reg[4][22]  ( .E(n5212), .D(\vrf/N40 ), .Q(
        \vrf/regTable[4][22] ) );
  LHQD1BWP \vrf/regTable_reg[4][23]  ( .E(n5212), .D(\vrf/N41 ), .Q(
        \vrf/regTable[4][23] ) );
  LHQD1BWP \vrf/regTable_reg[4][24]  ( .E(n5211), .D(\vrf/N42 ), .Q(
        \vrf/regTable[4][24] ) );
  LHQD1BWP \vrf/regTable_reg[4][25]  ( .E(n5211), .D(\vrf/N43 ), .Q(
        \vrf/regTable[4][25] ) );
  LHQD1BWP \vrf/regTable_reg[4][26]  ( .E(n5211), .D(\vrf/N44 ), .Q(
        \vrf/regTable[4][26] ) );
  LHQD1BWP \vrf/regTable_reg[4][27]  ( .E(n5211), .D(\vrf/N45 ), .Q(
        \vrf/regTable[4][27] ) );
  LHQD1BWP \vrf/regTable_reg[4][28]  ( .E(n5211), .D(\vrf/N46 ), .Q(
        \vrf/regTable[4][28] ) );
  LHQD1BWP \vrf/regTable_reg[4][29]  ( .E(n5211), .D(\vrf/N47 ), .Q(
        \vrf/regTable[4][29] ) );
  LHQD1BWP \vrf/regTable_reg[4][30]  ( .E(n5211), .D(\vrf/N48 ), .Q(
        \vrf/regTable[4][30] ) );
  LHQD1BWP \vrf/regTable_reg[4][31]  ( .E(n5211), .D(\vrf/N49 ), .Q(
        \vrf/regTable[4][31] ) );
  LHQD1BWP \vrf/regTable_reg[4][32]  ( .E(n5211), .D(\vrf/N50 ), .Q(
        \vrf/regTable[4][32] ) );
  LHQD1BWP \vrf/regTable_reg[4][33]  ( .E(n5211), .D(\vrf/N51 ), .Q(
        \vrf/regTable[4][33] ) );
  LHQD1BWP \vrf/regTable_reg[4][34]  ( .E(n5211), .D(\vrf/N52 ), .Q(
        \vrf/regTable[4][34] ) );
  LHQD1BWP \vrf/regTable_reg[4][35]  ( .E(n5210), .D(\vrf/N53 ), .Q(
        \vrf/regTable[4][35] ) );
  LHQD1BWP \vrf/regTable_reg[4][36]  ( .E(n5210), .D(\vrf/N54 ), .Q(
        \vrf/regTable[4][36] ) );
  LHQD1BWP \vrf/regTable_reg[4][37]  ( .E(n5210), .D(\vrf/N55 ), .Q(
        \vrf/regTable[4][37] ) );
  LHQD1BWP \vrf/regTable_reg[4][38]  ( .E(n5210), .D(\vrf/N56 ), .Q(
        \vrf/regTable[4][38] ) );
  LHQD1BWP \vrf/regTable_reg[4][39]  ( .E(n5210), .D(\vrf/N57 ), .Q(
        \vrf/regTable[4][39] ) );
  LHQD1BWP \vrf/regTable_reg[4][40]  ( .E(n5210), .D(\vrf/N58 ), .Q(
        \vrf/regTable[4][40] ) );
  LHQD1BWP \vrf/regTable_reg[4][41]  ( .E(n5210), .D(\vrf/N59 ), .Q(
        \vrf/regTable[4][41] ) );
  LHQD1BWP \vrf/regTable_reg[4][42]  ( .E(n5210), .D(\vrf/N60 ), .Q(
        \vrf/regTable[4][42] ) );
  LHQD1BWP \vrf/regTable_reg[4][43]  ( .E(n5210), .D(\vrf/N61 ), .Q(
        \vrf/regTable[4][43] ) );
  LHQD1BWP \vrf/regTable_reg[4][44]  ( .E(n5210), .D(\vrf/N62 ), .Q(
        \vrf/regTable[4][44] ) );
  LHQD1BWP \vrf/regTable_reg[4][45]  ( .E(n5210), .D(\vrf/N63 ), .Q(
        \vrf/regTable[4][45] ) );
  LHQD1BWP \vrf/regTable_reg[4][46]  ( .E(n5209), .D(\vrf/N64 ), .Q(
        \vrf/regTable[4][46] ) );
  LHQD1BWP \vrf/regTable_reg[4][47]  ( .E(n5209), .D(\vrf/N65 ), .Q(
        \vrf/regTable[4][47] ) );
  LHQD1BWP \vrf/regTable_reg[4][48]  ( .E(n5209), .D(\vrf/N66 ), .Q(
        \vrf/regTable[4][48] ) );
  LHQD1BWP \vrf/regTable_reg[4][49]  ( .E(n5209), .D(\vrf/N67 ), .Q(
        \vrf/regTable[4][49] ) );
  LHQD1BWP \vrf/regTable_reg[4][50]  ( .E(n5209), .D(\vrf/N68 ), .Q(
        \vrf/regTable[4][50] ) );
  LHQD1BWP \vrf/regTable_reg[4][51]  ( .E(n5209), .D(\vrf/N69 ), .Q(
        \vrf/regTable[4][51] ) );
  LHQD1BWP \vrf/regTable_reg[4][52]  ( .E(n5209), .D(\vrf/N70 ), .Q(
        \vrf/regTable[4][52] ) );
  LHQD1BWP \vrf/regTable_reg[4][53]  ( .E(n5209), .D(\vrf/N71 ), .Q(
        \vrf/regTable[4][53] ) );
  LHQD1BWP \vrf/regTable_reg[4][54]  ( .E(n5209), .D(\vrf/N72 ), .Q(
        \vrf/regTable[4][54] ) );
  LHQD1BWP \vrf/regTable_reg[4][55]  ( .E(n5209), .D(\vrf/N73 ), .Q(
        \vrf/regTable[4][55] ) );
  LHQD1BWP \vrf/regTable_reg[4][56]  ( .E(n5209), .D(\vrf/N74 ), .Q(
        \vrf/regTable[4][56] ) );
  LHQD1BWP \vrf/regTable_reg[4][57]  ( .E(n5208), .D(\vrf/N75 ), .Q(
        \vrf/regTable[4][57] ) );
  LHQD1BWP \vrf/regTable_reg[4][58]  ( .E(n5208), .D(\vrf/N76 ), .Q(
        \vrf/regTable[4][58] ) );
  LHQD1BWP \vrf/regTable_reg[4][59]  ( .E(n5208), .D(\vrf/N77 ), .Q(
        \vrf/regTable[4][59] ) );
  LHQD1BWP \vrf/regTable_reg[4][60]  ( .E(n5208), .D(\vrf/N78 ), .Q(
        \vrf/regTable[4][60] ) );
  LHQD1BWP \vrf/regTable_reg[4][61]  ( .E(n5208), .D(\vrf/N79 ), .Q(
        \vrf/regTable[4][61] ) );
  LHQD1BWP \vrf/regTable_reg[4][62]  ( .E(n5208), .D(\vrf/N80 ), .Q(
        \vrf/regTable[4][62] ) );
  LHQD1BWP \vrf/regTable_reg[4][63]  ( .E(n5208), .D(\vrf/N81 ), .Q(
        \vrf/regTable[4][63] ) );
  LHQD1BWP \vrf/regTable_reg[4][64]  ( .E(n5208), .D(\vrf/N82 ), .Q(
        \vrf/regTable[4][64] ) );
  LHQD1BWP \vrf/regTable_reg[4][65]  ( .E(n5208), .D(\vrf/N83 ), .Q(
        \vrf/regTable[4][65] ) );
  LHQD1BWP \vrf/regTable_reg[4][66]  ( .E(n5208), .D(\vrf/N84 ), .Q(
        \vrf/regTable[4][66] ) );
  LHQD1BWP \vrf/regTable_reg[4][67]  ( .E(n5208), .D(\vrf/N85 ), .Q(
        \vrf/regTable[4][67] ) );
  LHQD1BWP \vrf/regTable_reg[4][68]  ( .E(n5207), .D(\vrf/N86 ), .Q(
        \vrf/regTable[4][68] ) );
  LHQD1BWP \vrf/regTable_reg[4][69]  ( .E(n5207), .D(\vrf/N87 ), .Q(
        \vrf/regTable[4][69] ) );
  LHQD1BWP \vrf/regTable_reg[4][70]  ( .E(n5207), .D(\vrf/N88 ), .Q(
        \vrf/regTable[4][70] ) );
  LHQD1BWP \vrf/regTable_reg[4][71]  ( .E(n5207), .D(\vrf/N89 ), .Q(
        \vrf/regTable[4][71] ) );
  LHQD1BWP \vrf/regTable_reg[4][72]  ( .E(n5207), .D(\vrf/N90 ), .Q(
        \vrf/regTable[4][72] ) );
  LHQD1BWP \vrf/regTable_reg[4][73]  ( .E(n5207), .D(\vrf/N91 ), .Q(
        \vrf/regTable[4][73] ) );
  LHQD1BWP \vrf/regTable_reg[4][74]  ( .E(n5207), .D(\vrf/N92 ), .Q(
        \vrf/regTable[4][74] ) );
  LHQD1BWP \vrf/regTable_reg[4][75]  ( .E(n5207), .D(\vrf/N93 ), .Q(
        \vrf/regTable[4][75] ) );
  LHQD1BWP \vrf/regTable_reg[4][76]  ( .E(n5207), .D(\vrf/N94 ), .Q(
        \vrf/regTable[4][76] ) );
  LHQD1BWP \vrf/regTable_reg[4][77]  ( .E(n5207), .D(\vrf/N95 ), .Q(
        \vrf/regTable[4][77] ) );
  LHQD1BWP \vrf/regTable_reg[4][78]  ( .E(n5207), .D(\vrf/N96 ), .Q(
        \vrf/regTable[4][78] ) );
  LHQD1BWP \vrf/regTable_reg[4][79]  ( .E(n5206), .D(\vrf/N97 ), .Q(
        \vrf/regTable[4][79] ) );
  LHQD1BWP \vrf/regTable_reg[4][80]  ( .E(n5206), .D(\vrf/N98 ), .Q(
        \vrf/regTable[4][80] ) );
  LHQD1BWP \vrf/regTable_reg[4][81]  ( .E(n5206), .D(\vrf/N99 ), .Q(
        \vrf/regTable[4][81] ) );
  LHQD1BWP \vrf/regTable_reg[4][82]  ( .E(n5206), .D(\vrf/N100 ), .Q(
        \vrf/regTable[4][82] ) );
  LHQD1BWP \vrf/regTable_reg[4][83]  ( .E(n5206), .D(\vrf/N101 ), .Q(
        \vrf/regTable[4][83] ) );
  LHQD1BWP \vrf/regTable_reg[4][84]  ( .E(n5206), .D(\vrf/N102 ), .Q(
        \vrf/regTable[4][84] ) );
  LHQD1BWP \vrf/regTable_reg[4][85]  ( .E(n5206), .D(\vrf/N103 ), .Q(
        \vrf/regTable[4][85] ) );
  LHQD1BWP \vrf/regTable_reg[4][86]  ( .E(n5206), .D(\vrf/N104 ), .Q(
        \vrf/regTable[4][86] ) );
  LHQD1BWP \vrf/regTable_reg[4][87]  ( .E(n5206), .D(\vrf/N105 ), .Q(
        \vrf/regTable[4][87] ) );
  LHQD1BWP \vrf/regTable_reg[4][88]  ( .E(n5206), .D(\vrf/N106 ), .Q(
        \vrf/regTable[4][88] ) );
  LHQD1BWP \vrf/regTable_reg[4][89]  ( .E(n5206), .D(\vrf/N107 ), .Q(
        \vrf/regTable[4][89] ) );
  LHQD1BWP \vrf/regTable_reg[4][90]  ( .E(n5205), .D(\vrf/N108 ), .Q(
        \vrf/regTable[4][90] ) );
  LHQD1BWP \vrf/regTable_reg[4][91]  ( .E(n5205), .D(\vrf/N109 ), .Q(
        \vrf/regTable[4][91] ) );
  LHQD1BWP \vrf/regTable_reg[4][92]  ( .E(n5205), .D(\vrf/N110 ), .Q(
        \vrf/regTable[4][92] ) );
  LHQD1BWP \vrf/regTable_reg[4][93]  ( .E(n5205), .D(\vrf/N111 ), .Q(
        \vrf/regTable[4][93] ) );
  LHQD1BWP \vrf/regTable_reg[4][94]  ( .E(n5205), .D(\vrf/N112 ), .Q(
        \vrf/regTable[4][94] ) );
  LHQD1BWP \vrf/regTable_reg[4][95]  ( .E(n5205), .D(\vrf/N113 ), .Q(
        \vrf/regTable[4][95] ) );
  LHQD1BWP \vrf/regTable_reg[4][96]  ( .E(n5205), .D(\vrf/N114 ), .Q(
        \vrf/regTable[4][96] ) );
  LHQD1BWP \vrf/regTable_reg[4][97]  ( .E(n5205), .D(\vrf/N115 ), .Q(
        \vrf/regTable[4][97] ) );
  LHQD1BWP \vrf/regTable_reg[4][98]  ( .E(n5205), .D(\vrf/N116 ), .Q(
        \vrf/regTable[4][98] ) );
  LHQD1BWP \vrf/regTable_reg[4][99]  ( .E(n5205), .D(\vrf/N118 ), .Q(
        \vrf/regTable[4][99] ) );
  LHQD1BWP \vrf/regTable_reg[4][100]  ( .E(n5215), .D(\vrf/N119 ), .Q(
        \vrf/regTable[4][100] ) );
  LHQD1BWP \vrf/regTable_reg[4][101]  ( .E(n5215), .D(\vrf/N120 ), .Q(
        \vrf/regTable[4][101] ) );
  LHQD1BWP \vrf/regTable_reg[4][102]  ( .E(n5215), .D(\vrf/N121 ), .Q(
        \vrf/regTable[4][102] ) );
  LHQD1BWP \vrf/regTable_reg[4][103]  ( .E(n5215), .D(\vrf/N122 ), .Q(
        \vrf/regTable[4][103] ) );
  LHQD1BWP \vrf/regTable_reg[4][104]  ( .E(n5215), .D(\vrf/N123 ), .Q(
        \vrf/regTable[4][104] ) );
  LHQD1BWP \vrf/regTable_reg[4][105]  ( .E(n5214), .D(\vrf/N124 ), .Q(
        \vrf/regTable[4][105] ) );
  LHQD1BWP \vrf/regTable_reg[4][106]  ( .E(n5214), .D(\vrf/N125 ), .Q(
        \vrf/regTable[4][106] ) );
  LHQD1BWP \vrf/regTable_reg[4][107]  ( .E(n5214), .D(\vrf/N126 ), .Q(
        \vrf/regTable[4][107] ) );
  LHQD1BWP \vrf/regTable_reg[4][108]  ( .E(n5214), .D(\vrf/N127 ), .Q(
        \vrf/regTable[4][108] ) );
  LHQD1BWP \vrf/regTable_reg[4][109]  ( .E(n5214), .D(\vrf/N128 ), .Q(
        \vrf/regTable[4][109] ) );
  LHQD1BWP \vrf/regTable_reg[4][110]  ( .E(n5214), .D(\vrf/N129 ), .Q(
        \vrf/regTable[4][110] ) );
  LHQD1BWP \vrf/regTable_reg[4][111]  ( .E(n5214), .D(\vrf/N130 ), .Q(
        \vrf/regTable[4][111] ) );
  LHQD1BWP \vrf/regTable_reg[4][112]  ( .E(n5214), .D(\vrf/N131 ), .Q(
        \vrf/regTable[4][112] ) );
  LHQD1BWP \vrf/regTable_reg[4][113]  ( .E(n5214), .D(\vrf/N132 ), .Q(
        \vrf/regTable[4][113] ) );
  LHQD1BWP \vrf/regTable_reg[4][114]  ( .E(n5214), .D(\vrf/N133 ), .Q(
        \vrf/regTable[4][114] ) );
  LHQD1BWP \vrf/regTable_reg[4][115]  ( .E(n5214), .D(\vrf/N134 ), .Q(
        \vrf/regTable[4][115] ) );
  LHQD1BWP \vrf/regTable_reg[4][116]  ( .E(n5213), .D(\vrf/N135 ), .Q(
        \vrf/regTable[4][116] ) );
  LHQD1BWP \vrf/regTable_reg[4][117]  ( .E(n5213), .D(\vrf/N136 ), .Q(
        \vrf/regTable[4][117] ) );
  LHQD1BWP \vrf/regTable_reg[4][118]  ( .E(n5213), .D(\vrf/N137 ), .Q(
        \vrf/regTable[4][118] ) );
  LHQD1BWP \vrf/regTable_reg[4][119]  ( .E(n5213), .D(\vrf/N138 ), .Q(
        \vrf/regTable[4][119] ) );
  LHQD1BWP \vrf/regTable_reg[4][120]  ( .E(n5213), .D(\vrf/N139 ), .Q(
        \vrf/regTable[4][120] ) );
  LHQD1BWP \vrf/regTable_reg[4][121]  ( .E(n5213), .D(\vrf/N140 ), .Q(
        \vrf/regTable[4][121] ) );
  LHQD1BWP \vrf/regTable_reg[4][122]  ( .E(n5213), .D(\vrf/N141 ), .Q(
        \vrf/regTable[4][122] ) );
  LHQD1BWP \vrf/regTable_reg[4][123]  ( .E(n5213), .D(\vrf/N142 ), .Q(
        \vrf/regTable[4][123] ) );
  LHQD1BWP \vrf/regTable_reg[4][124]  ( .E(n5213), .D(\vrf/N143 ), .Q(
        \vrf/regTable[4][124] ) );
  LHQD1BWP \vrf/regTable_reg[4][125]  ( .E(n5213), .D(\vrf/N144 ), .Q(
        \vrf/regTable[4][125] ) );
  LHQD1BWP \vrf/regTable_reg[4][126]  ( .E(n5213), .D(\vrf/N145 ), .Q(
        \vrf/regTable[4][126] ) );
  LHQD1BWP \vrf/regTable_reg[4][127]  ( .E(n5212), .D(\vrf/N146 ), .Q(
        \vrf/regTable[4][127] ) );
  LHQD1BWP \vrf/regTable_reg[4][128]  ( .E(n5215), .D(\vrf/N147 ), .Q(
        \vrf/regTable[4][128] ) );
  LHQD1BWP \vrf/regTable_reg[4][129]  ( .E(n5215), .D(\vrf/N148 ), .Q(
        \vrf/regTable[4][129] ) );
  LHQD1BWP \vrf/regTable_reg[4][130]  ( .E(n5215), .D(\vrf/N149 ), .Q(
        \vrf/regTable[4][130] ) );
  LHQD1BWP \vrf/regTable_reg[4][131]  ( .E(n5215), .D(\vrf/N150 ), .Q(
        \vrf/regTable[4][131] ) );
  LHQD1BWP \vrf/regTable_reg[4][132]  ( .E(n5215), .D(\vrf/N151 ), .Q(
        \vrf/regTable[4][132] ) );
  LHQD1BWP \vrf/regTable_reg[4][133]  ( .E(n5215), .D(\vrf/N152 ), .Q(
        \vrf/regTable[4][133] ) );
  LHQD1BWP \vrf/regTable_reg[4][134]  ( .E(n5216), .D(\vrf/N153 ), .Q(
        \vrf/regTable[4][134] ) );
  LHQD1BWP \vrf/regTable_reg[4][135]  ( .E(n5216), .D(\vrf/N154 ), .Q(
        \vrf/regTable[4][135] ) );
  LHQD1BWP \vrf/regTable_reg[4][136]  ( .E(n5216), .D(\vrf/N155 ), .Q(
        \vrf/regTable[4][136] ) );
  LHQD1BWP \vrf/regTable_reg[4][137]  ( .E(n5216), .D(\vrf/N156 ), .Q(
        \vrf/regTable[4][137] ) );
  LHQD1BWP \vrf/regTable_reg[4][138]  ( .E(n5216), .D(\vrf/N157 ), .Q(
        \vrf/regTable[4][138] ) );
  LHQD1BWP \vrf/regTable_reg[4][139]  ( .E(n5216), .D(\vrf/N158 ), .Q(
        \vrf/regTable[4][139] ) );
  LHQD1BWP \vrf/regTable_reg[4][140]  ( .E(n5216), .D(\vrf/N159 ), .Q(
        \vrf/regTable[4][140] ) );
  LHQD1BWP \vrf/regTable_reg[4][141]  ( .E(n5216), .D(\vrf/N160 ), .Q(
        \vrf/regTable[4][141] ) );
  LHQD1BWP \vrf/regTable_reg[4][142]  ( .E(n5216), .D(\vrf/N161 ), .Q(
        \vrf/regTable[4][142] ) );
  LHQD1BWP \vrf/regTable_reg[4][143]  ( .E(n5216), .D(\vrf/N162 ), .Q(
        \vrf/regTable[4][143] ) );
  LHQD1BWP \vrf/regTable_reg[4][144]  ( .E(n5216), .D(\vrf/N163 ), .Q(
        \vrf/regTable[4][144] ) );
  LHQD1BWP \vrf/regTable_reg[4][145]  ( .E(n5216), .D(\vrf/N164 ), .Q(
        \vrf/regTable[4][145] ) );
  LHQD1BWP \vrf/regTable_reg[4][146]  ( .E(n5217), .D(\vrf/N165 ), .Q(
        \vrf/regTable[4][146] ) );
  LHQD1BWP \vrf/regTable_reg[4][147]  ( .E(n5217), .D(\vrf/N166 ), .Q(
        \vrf/regTable[4][147] ) );
  LHQD1BWP \vrf/regTable_reg[4][148]  ( .E(n5217), .D(\vrf/N167 ), .Q(
        \vrf/regTable[4][148] ) );
  LHQD1BWP \vrf/regTable_reg[4][149]  ( .E(n5217), .D(\vrf/N168 ), .Q(
        \vrf/regTable[4][149] ) );
  LHQD1BWP \vrf/regTable_reg[4][150]  ( .E(n5217), .D(\vrf/N169 ), .Q(
        \vrf/regTable[4][150] ) );
  LHQD1BWP \vrf/regTable_reg[4][151]  ( .E(n5217), .D(\vrf/N170 ), .Q(
        \vrf/regTable[4][151] ) );
  LHQD1BWP \vrf/regTable_reg[4][152]  ( .E(n5217), .D(\vrf/N171 ), .Q(
        \vrf/regTable[4][152] ) );
  LHQD1BWP \vrf/regTable_reg[4][153]  ( .E(n5217), .D(\vrf/N172 ), .Q(
        \vrf/regTable[4][153] ) );
  LHQD1BWP \vrf/regTable_reg[4][154]  ( .E(n5217), .D(\vrf/N173 ), .Q(
        \vrf/regTable[4][154] ) );
  LHQD1BWP \vrf/regTable_reg[4][155]  ( .E(n5217), .D(\vrf/N174 ), .Q(
        \vrf/regTable[4][155] ) );
  LHQD1BWP \vrf/regTable_reg[4][156]  ( .E(n5217), .D(\vrf/N175 ), .Q(
        \vrf/regTable[4][156] ) );
  LHQD1BWP \vrf/regTable_reg[4][157]  ( .E(n5217), .D(\vrf/N176 ), .Q(
        \vrf/regTable[4][157] ) );
  LHQD1BWP \vrf/regTable_reg[4][158]  ( .E(n5218), .D(\vrf/N177 ), .Q(
        \vrf/regTable[4][158] ) );
  LHQD1BWP \vrf/regTable_reg[4][159]  ( .E(n5218), .D(\vrf/N178 ), .Q(
        \vrf/regTable[4][159] ) );
  LHQD1BWP \vrf/regTable_reg[4][160]  ( .E(n5218), .D(\vrf/N179 ), .Q(
        \vrf/regTable[4][160] ) );
  LHQD1BWP \vrf/regTable_reg[4][161]  ( .E(n5218), .D(\vrf/N180 ), .Q(
        \vrf/regTable[4][161] ) );
  LHQD1BWP \vrf/regTable_reg[4][162]  ( .E(n5218), .D(\vrf/N181 ), .Q(
        \vrf/regTable[4][162] ) );
  LHQD1BWP \vrf/regTable_reg[4][163]  ( .E(n5218), .D(\vrf/N182 ), .Q(
        \vrf/regTable[4][163] ) );
  LHQD1BWP \vrf/regTable_reg[4][164]  ( .E(n5218), .D(\vrf/N183 ), .Q(
        \vrf/regTable[4][164] ) );
  LHQD1BWP \vrf/regTable_reg[4][165]  ( .E(n5218), .D(\vrf/N184 ), .Q(
        \vrf/regTable[4][165] ) );
  LHQD1BWP \vrf/regTable_reg[4][166]  ( .E(n5218), .D(\vrf/N185 ), .Q(
        \vrf/regTable[4][166] ) );
  LHQD1BWP \vrf/regTable_reg[4][167]  ( .E(n5218), .D(\vrf/N186 ), .Q(
        \vrf/regTable[4][167] ) );
  LHQD1BWP \vrf/regTable_reg[4][168]  ( .E(n5218), .D(\vrf/N187 ), .Q(
        \vrf/regTable[4][168] ) );
  LHQD1BWP \vrf/regTable_reg[4][169]  ( .E(n5218), .D(\vrf/N188 ), .Q(
        \vrf/regTable[4][169] ) );
  LHQD1BWP \vrf/regTable_reg[4][170]  ( .E(n5219), .D(\vrf/N189 ), .Q(
        \vrf/regTable[4][170] ) );
  LHQD1BWP \vrf/regTable_reg[4][171]  ( .E(n5219), .D(\vrf/N190 ), .Q(
        \vrf/regTable[4][171] ) );
  LHQD1BWP \vrf/regTable_reg[4][172]  ( .E(n5219), .D(\vrf/N191 ), .Q(
        \vrf/regTable[4][172] ) );
  LHQD1BWP \vrf/regTable_reg[4][173]  ( .E(n5219), .D(\vrf/N192 ), .Q(
        \vrf/regTable[4][173] ) );
  LHQD1BWP \vrf/regTable_reg[4][174]  ( .E(n5219), .D(\vrf/N193 ), .Q(
        \vrf/regTable[4][174] ) );
  LHQD1BWP \vrf/regTable_reg[4][175]  ( .E(n5219), .D(\vrf/N194 ), .Q(
        \vrf/regTable[4][175] ) );
  LHQD1BWP \vrf/regTable_reg[4][176]  ( .E(n5219), .D(\vrf/N195 ), .Q(
        \vrf/regTable[4][176] ) );
  LHQD1BWP \vrf/regTable_reg[4][177]  ( .E(n5219), .D(\vrf/N196 ), .Q(
        \vrf/regTable[4][177] ) );
  LHQD1BWP \vrf/regTable_reg[4][178]  ( .E(n5219), .D(\vrf/N197 ), .Q(
        \vrf/regTable[4][178] ) );
  LHQD1BWP \vrf/regTable_reg[4][179]  ( .E(n5219), .D(\vrf/N198 ), .Q(
        \vrf/regTable[4][179] ) );
  LHQD1BWP \vrf/regTable_reg[4][180]  ( .E(n5219), .D(\vrf/N199 ), .Q(
        \vrf/regTable[4][180] ) );
  LHQD1BWP \vrf/regTable_reg[4][181]  ( .E(n5219), .D(\vrf/N200 ), .Q(
        \vrf/regTable[4][181] ) );
  LHQD1BWP \vrf/regTable_reg[4][182]  ( .E(n5220), .D(\vrf/N201 ), .Q(
        \vrf/regTable[4][182] ) );
  LHQD1BWP \vrf/regTable_reg[4][183]  ( .E(n5220), .D(\vrf/N202 ), .Q(
        \vrf/regTable[4][183] ) );
  LHQD1BWP \vrf/regTable_reg[4][184]  ( .E(n5220), .D(\vrf/N203 ), .Q(
        \vrf/regTable[4][184] ) );
  LHQD1BWP \vrf/regTable_reg[4][185]  ( .E(n5220), .D(\vrf/N204 ), .Q(
        \vrf/regTable[4][185] ) );
  LHQD1BWP \vrf/regTable_reg[4][186]  ( .E(n5220), .D(\vrf/N205 ), .Q(
        \vrf/regTable[4][186] ) );
  LHQD1BWP \vrf/regTable_reg[4][187]  ( .E(n5220), .D(\vrf/N206 ), .Q(
        \vrf/regTable[4][187] ) );
  LHQD1BWP \vrf/regTable_reg[4][188]  ( .E(n5220), .D(\vrf/N207 ), .Q(
        \vrf/regTable[4][188] ) );
  LHQD1BWP \vrf/regTable_reg[4][189]  ( .E(n5220), .D(\vrf/N208 ), .Q(
        \vrf/regTable[4][189] ) );
  LHQD1BWP \vrf/regTable_reg[4][190]  ( .E(n5220), .D(\vrf/N209 ), .Q(
        \vrf/regTable[4][190] ) );
  LHQD1BWP \vrf/regTable_reg[4][191]  ( .E(n5220), .D(\vrf/N210 ), .Q(
        \vrf/regTable[4][191] ) );
  LHQD1BWP \vrf/regTable_reg[4][192]  ( .E(n5220), .D(\vrf/N211 ), .Q(
        \vrf/regTable[4][192] ) );
  LHQD1BWP \vrf/regTable_reg[4][193]  ( .E(n5220), .D(\vrf/N212 ), .Q(
        \vrf/regTable[4][193] ) );
  LHQD1BWP \vrf/regTable_reg[4][194]  ( .E(n5221), .D(\vrf/N213 ), .Q(
        \vrf/regTable[4][194] ) );
  LHQD1BWP \vrf/regTable_reg[4][195]  ( .E(n5221), .D(\vrf/N214 ), .Q(
        \vrf/regTable[4][195] ) );
  LHQD1BWP \vrf/regTable_reg[4][196]  ( .E(n5221), .D(\vrf/N215 ), .Q(
        \vrf/regTable[4][196] ) );
  LHQD1BWP \vrf/regTable_reg[4][197]  ( .E(n5221), .D(\vrf/N216 ), .Q(
        \vrf/regTable[4][197] ) );
  LHQD1BWP \vrf/regTable_reg[4][198]  ( .E(n5221), .D(\vrf/N218 ), .Q(
        \vrf/regTable[4][198] ) );
  LHQD1BWP \vrf/regTable_reg[4][199]  ( .E(n5221), .D(\vrf/N219 ), .Q(
        \vrf/regTable[4][199] ) );
  LHQD1BWP \vrf/regTable_reg[4][200]  ( .E(n5221), .D(\vrf/N220 ), .Q(
        \vrf/regTable[4][200] ) );
  LHQD1BWP \vrf/regTable_reg[4][201]  ( .E(n5221), .D(\vrf/N221 ), .Q(
        \vrf/regTable[4][201] ) );
  LHQD1BWP \vrf/regTable_reg[4][202]  ( .E(n5221), .D(\vrf/N222 ), .Q(
        \vrf/regTable[4][202] ) );
  LHQD1BWP \vrf/regTable_reg[4][203]  ( .E(n5221), .D(\vrf/N223 ), .Q(
        \vrf/regTable[4][203] ) );
  LHQD1BWP \vrf/regTable_reg[4][204]  ( .E(n5221), .D(\vrf/N224 ), .Q(
        \vrf/regTable[4][204] ) );
  LHQD1BWP \vrf/regTable_reg[4][205]  ( .E(n5221), .D(\vrf/N225 ), .Q(
        \vrf/regTable[4][205] ) );
  LHQD1BWP \vrf/regTable_reg[4][206]  ( .E(n5222), .D(\vrf/N226 ), .Q(
        \vrf/regTable[4][206] ) );
  LHQD1BWP \vrf/regTable_reg[4][207]  ( .E(n5222), .D(\vrf/N227 ), .Q(
        \vrf/regTable[4][207] ) );
  LHQD1BWP \vrf/regTable_reg[4][208]  ( .E(n5222), .D(\vrf/N228 ), .Q(
        \vrf/regTable[4][208] ) );
  LHQD1BWP \vrf/regTable_reg[4][209]  ( .E(n5222), .D(\vrf/N229 ), .Q(
        \vrf/regTable[4][209] ) );
  LHQD1BWP \vrf/regTable_reg[4][210]  ( .E(n5222), .D(\vrf/N230 ), .Q(
        \vrf/regTable[4][210] ) );
  LHQD1BWP \vrf/regTable_reg[4][211]  ( .E(n5222), .D(\vrf/N231 ), .Q(
        \vrf/regTable[4][211] ) );
  LHQD1BWP \vrf/regTable_reg[4][212]  ( .E(n5222), .D(\vrf/N232 ), .Q(
        \vrf/regTable[4][212] ) );
  LHQD1BWP \vrf/regTable_reg[4][213]  ( .E(n5222), .D(\vrf/N233 ), .Q(
        \vrf/regTable[4][213] ) );
  LHQD1BWP \vrf/regTable_reg[4][214]  ( .E(n5222), .D(\vrf/N234 ), .Q(
        \vrf/regTable[4][214] ) );
  LHQD1BWP \vrf/regTable_reg[4][215]  ( .E(n5222), .D(\vrf/N235 ), .Q(
        \vrf/regTable[4][215] ) );
  LHQD1BWP \vrf/regTable_reg[4][216]  ( .E(n5222), .D(\vrf/N236 ), .Q(
        \vrf/regTable[4][216] ) );
  LHQD1BWP \vrf/regTable_reg[4][217]  ( .E(n5222), .D(\vrf/N237 ), .Q(
        \vrf/regTable[4][217] ) );
  LHQD1BWP \vrf/regTable_reg[4][218]  ( .E(n5223), .D(\vrf/N238 ), .Q(
        \vrf/regTable[4][218] ) );
  LHQD1BWP \vrf/regTable_reg[4][219]  ( .E(n5223), .D(\vrf/N239 ), .Q(
        \vrf/regTable[4][219] ) );
  LHQD1BWP \vrf/regTable_reg[4][220]  ( .E(n5223), .D(\vrf/N240 ), .Q(
        \vrf/regTable[4][220] ) );
  LHQD1BWP \vrf/regTable_reg[4][221]  ( .E(n5223), .D(\vrf/N241 ), .Q(
        \vrf/regTable[4][221] ) );
  LHQD1BWP \vrf/regTable_reg[4][222]  ( .E(n5223), .D(\vrf/N242 ), .Q(
        \vrf/regTable[4][222] ) );
  LHQD1BWP \vrf/regTable_reg[4][223]  ( .E(n5223), .D(\vrf/N243 ), .Q(
        \vrf/regTable[4][223] ) );
  LHQD1BWP \vrf/regTable_reg[4][224]  ( .E(n5223), .D(\vrf/N244 ), .Q(
        \vrf/regTable[4][224] ) );
  LHQD1BWP \vrf/regTable_reg[4][225]  ( .E(n5223), .D(\vrf/N245 ), .Q(
        \vrf/regTable[4][225] ) );
  LHQD1BWP \vrf/regTable_reg[4][226]  ( .E(n5223), .D(\vrf/N246 ), .Q(
        \vrf/regTable[4][226] ) );
  LHQD1BWP \vrf/regTable_reg[4][227]  ( .E(n5223), .D(\vrf/N247 ), .Q(
        \vrf/regTable[4][227] ) );
  LHQD1BWP \vrf/regTable_reg[4][228]  ( .E(n5223), .D(\vrf/N248 ), .Q(
        \vrf/regTable[4][228] ) );
  LHQD1BWP \vrf/regTable_reg[4][229]  ( .E(n5223), .D(\vrf/N249 ), .Q(
        \vrf/regTable[4][229] ) );
  LHQD1BWP \vrf/regTable_reg[4][230]  ( .E(n5224), .D(\vrf/N250 ), .Q(
        \vrf/regTable[4][230] ) );
  LHQD1BWP \vrf/regTable_reg[4][231]  ( .E(n5224), .D(\vrf/N251 ), .Q(
        \vrf/regTable[4][231] ) );
  LHQD1BWP \vrf/regTable_reg[4][232]  ( .E(n5224), .D(\vrf/N252 ), .Q(
        \vrf/regTable[4][232] ) );
  LHQD1BWP \vrf/regTable_reg[4][233]  ( .E(n5224), .D(\vrf/N253 ), .Q(
        \vrf/regTable[4][233] ) );
  LHQD1BWP \vrf/regTable_reg[4][234]  ( .E(n5224), .D(\vrf/N254 ), .Q(
        \vrf/regTable[4][234] ) );
  LHQD1BWP \vrf/regTable_reg[4][235]  ( .E(n5224), .D(\vrf/N255 ), .Q(
        \vrf/regTable[4][235] ) );
  LHQD1BWP \vrf/regTable_reg[4][236]  ( .E(n5224), .D(\vrf/N256 ), .Q(
        \vrf/regTable[4][236] ) );
  LHQD1BWP \vrf/regTable_reg[4][237]  ( .E(n5224), .D(\vrf/N257 ), .Q(
        \vrf/regTable[4][237] ) );
  LHQD1BWP \vrf/regTable_reg[4][238]  ( .E(n5224), .D(\vrf/N258 ), .Q(
        \vrf/regTable[4][238] ) );
  LHQD1BWP \vrf/regTable_reg[4][239]  ( .E(n5224), .D(\vrf/N259 ), .Q(
        \vrf/regTable[4][239] ) );
  LHQD1BWP \vrf/regTable_reg[4][240]  ( .E(n5224), .D(\vrf/N260 ), .Q(
        \vrf/regTable[4][240] ) );
  LHQD1BWP \vrf/regTable_reg[4][241]  ( .E(n5224), .D(\vrf/N261 ), .Q(
        \vrf/regTable[4][241] ) );
  LHQD1BWP \vrf/regTable_reg[4][242]  ( .E(n5225), .D(\vrf/N262 ), .Q(
        \vrf/regTable[4][242] ) );
  LHQD1BWP \vrf/regTable_reg[4][243]  ( .E(n5225), .D(\vrf/N263 ), .Q(
        \vrf/regTable[4][243] ) );
  LHQD1BWP \vrf/regTable_reg[4][244]  ( .E(n5225), .D(\vrf/N264 ), .Q(
        \vrf/regTable[4][244] ) );
  LHQD1BWP \vrf/regTable_reg[4][245]  ( .E(n5225), .D(\vrf/N265 ), .Q(
        \vrf/regTable[4][245] ) );
  LHQD1BWP \vrf/regTable_reg[4][246]  ( .E(n5225), .D(\vrf/N266 ), .Q(
        \vrf/regTable[4][246] ) );
  LHQD1BWP \vrf/regTable_reg[4][247]  ( .E(n5225), .D(\vrf/N267 ), .Q(
        \vrf/regTable[4][247] ) );
  LHQD1BWP \vrf/regTable_reg[4][248]  ( .E(n5225), .D(\vrf/N268 ), .Q(
        \vrf/regTable[4][248] ) );
  LHQD1BWP \vrf/regTable_reg[4][249]  ( .E(n5225), .D(\vrf/N269 ), .Q(
        \vrf/regTable[4][249] ) );
  LHQD1BWP \vrf/regTable_reg[4][250]  ( .E(n5225), .D(\vrf/N270 ), .Q(
        \vrf/regTable[4][250] ) );
  LHQD1BWP \vrf/regTable_reg[4][251]  ( .E(n5225), .D(\vrf/N271 ), .Q(
        \vrf/regTable[4][251] ) );
  LHQD1BWP \vrf/regTable_reg[4][252]  ( .E(n5225), .D(\vrf/N272 ), .Q(
        \vrf/regTable[4][252] ) );
  LHQD1BWP \vrf/regTable_reg[4][253]  ( .E(n5225), .D(\vrf/N273 ), .Q(
        \vrf/regTable[4][253] ) );
  LHQD1BWP \vrf/regTable_reg[0][0]  ( .E(n5351), .D(\vrf/N18 ), .Q(
        \vrf/regTable[0][0] ) );
  LHQD1BWP \vrf/regTable_reg[0][1]  ( .E(n5348), .D(\vrf/N19 ), .Q(
        \vrf/regTable[0][1] ) );
  LHQD1BWP \vrf/regTable_reg[0][2]  ( .E(n5347), .D(\vrf/N20 ), .Q(
        \vrf/regTable[0][2] ) );
  LHQD1BWP \vrf/regTable_reg[0][3]  ( .E(n5346), .D(\vrf/N21 ), .Q(
        \vrf/regTable[0][3] ) );
  LHQD1BWP \vrf/regTable_reg[0][4]  ( .E(n5345), .D(\vrf/N22 ), .Q(
        \vrf/regTable[0][4] ) );
  LHQD1BWP \vrf/regTable_reg[0][5]  ( .E(n5344), .D(\vrf/N23 ), .Q(
        \vrf/regTable[0][5] ) );
  LHQD1BWP \vrf/regTable_reg[0][6]  ( .E(n5343), .D(\vrf/N24 ), .Q(
        \vrf/regTable[0][6] ) );
  LHQD1BWP \vrf/regTable_reg[0][7]  ( .E(n5342), .D(\vrf/N25 ), .Q(
        \vrf/regTable[0][7] ) );
  LHQD1BWP \vrf/regTable_reg[0][8]  ( .E(n5341), .D(\vrf/N26 ), .Q(
        \vrf/regTable[0][8] ) );
  LHQD1BWP \vrf/regTable_reg[0][9]  ( .E(n5341), .D(\vrf/N27 ), .Q(
        \vrf/regTable[0][9] ) );
  LHQD1BWP \vrf/regTable_reg[0][10]  ( .E(n5350), .D(\vrf/N28 ), .Q(
        \vrf/regTable[0][10] ) );
  LHQD1BWP \vrf/regTable_reg[0][11]  ( .E(n5349), .D(\vrf/N29 ), .Q(
        \vrf/regTable[0][11] ) );
  LHQD1BWP \vrf/regTable_reg[0][12]  ( .E(n5348), .D(\vrf/N30 ), .Q(
        \vrf/regTable[0][12] ) );
  LHQD1BWP \vrf/regTable_reg[0][13]  ( .E(n5348), .D(\vrf/N31 ), .Q(
        \vrf/regTable[0][13] ) );
  LHQD1BWP \vrf/regTable_reg[0][14]  ( .E(n5348), .D(\vrf/N32 ), .Q(
        \vrf/regTable[0][14] ) );
  LHQD1BWP \vrf/regTable_reg[0][17]  ( .E(n5348), .D(\vrf/N35 ), .Q(
        \vrf/regTable[0][17] ) );
  LHQD1BWP \vrf/regTable_reg[0][18]  ( .E(n5348), .D(\vrf/N36 ), .Q(
        \vrf/regTable[0][18] ) );
  LHQD1BWP \vrf/regTable_reg[0][19]  ( .E(n5348), .D(\vrf/N37 ), .Q(
        \vrf/regTable[0][19] ) );
  LHQD1BWP \vrf/regTable_reg[0][20]  ( .E(n5348), .D(\vrf/N38 ), .Q(
        \vrf/regTable[0][20] ) );
  LHQD1BWP \vrf/regTable_reg[0][21]  ( .E(n5348), .D(\vrf/N39 ), .Q(
        \vrf/regTable[0][21] ) );
  LHQD1BWP \vrf/regTable_reg[0][22]  ( .E(n5348), .D(\vrf/N40 ), .Q(
        \vrf/regTable[0][22] ) );
  LHQD1BWP \vrf/regTable_reg[0][23]  ( .E(n5348), .D(\vrf/N41 ), .Q(
        \vrf/regTable[0][23] ) );
  LHQD1BWP \vrf/regTable_reg[0][24]  ( .E(n5347), .D(\vrf/N42 ), .Q(
        \vrf/regTable[0][24] ) );
  LHQD1BWP \vrf/regTable_reg[0][25]  ( .E(n5347), .D(\vrf/N43 ), .Q(
        \vrf/regTable[0][25] ) );
  LHQD1BWP \vrf/regTable_reg[0][26]  ( .E(n5347), .D(\vrf/N44 ), .Q(
        \vrf/regTable[0][26] ) );
  LHQD1BWP \vrf/regTable_reg[0][27]  ( .E(n5347), .D(\vrf/N45 ), .Q(
        \vrf/regTable[0][27] ) );
  LHQD1BWP \vrf/regTable_reg[0][28]  ( .E(n5347), .D(\vrf/N46 ), .Q(
        \vrf/regTable[0][28] ) );
  LHQD1BWP \vrf/regTable_reg[0][29]  ( .E(n5347), .D(\vrf/N47 ), .Q(
        \vrf/regTable[0][29] ) );
  LHQD1BWP \vrf/regTable_reg[0][30]  ( .E(n5347), .D(\vrf/N48 ), .Q(
        \vrf/regTable[0][30] ) );
  LHQD1BWP \vrf/regTable_reg[0][31]  ( .E(n5347), .D(\vrf/N49 ), .Q(
        \vrf/regTable[0][31] ) );
  LHQD1BWP \vrf/regTable_reg[0][32]  ( .E(n5347), .D(\vrf/N50 ), .Q(
        \vrf/regTable[0][32] ) );
  LHQD1BWP \vrf/regTable_reg[0][33]  ( .E(n5347), .D(\vrf/N51 ), .Q(
        \vrf/regTable[0][33] ) );
  LHQD1BWP \vrf/regTable_reg[0][34]  ( .E(n5347), .D(\vrf/N52 ), .Q(
        \vrf/regTable[0][34] ) );
  LHQD1BWP \vrf/regTable_reg[0][35]  ( .E(n5346), .D(\vrf/N53 ), .Q(
        \vrf/regTable[0][35] ) );
  LHQD1BWP \vrf/regTable_reg[0][36]  ( .E(n5346), .D(\vrf/N54 ), .Q(
        \vrf/regTable[0][36] ) );
  LHQD1BWP \vrf/regTable_reg[0][37]  ( .E(n5346), .D(\vrf/N55 ), .Q(
        \vrf/regTable[0][37] ) );
  LHQD1BWP \vrf/regTable_reg[0][38]  ( .E(n5346), .D(\vrf/N56 ), .Q(
        \vrf/regTable[0][38] ) );
  LHQD1BWP \vrf/regTable_reg[0][39]  ( .E(n5346), .D(\vrf/N57 ), .Q(
        \vrf/regTable[0][39] ) );
  LHQD1BWP \vrf/regTable_reg[0][40]  ( .E(n5346), .D(\vrf/N58 ), .Q(
        \vrf/regTable[0][40] ) );
  LHQD1BWP \vrf/regTable_reg[0][41]  ( .E(n5346), .D(\vrf/N59 ), .Q(
        \vrf/regTable[0][41] ) );
  LHQD1BWP \vrf/regTable_reg[0][42]  ( .E(n5346), .D(\vrf/N60 ), .Q(
        \vrf/regTable[0][42] ) );
  LHQD1BWP \vrf/regTable_reg[0][43]  ( .E(n5346), .D(\vrf/N61 ), .Q(
        \vrf/regTable[0][43] ) );
  LHQD1BWP \vrf/regTable_reg[0][44]  ( .E(n5346), .D(\vrf/N62 ), .Q(
        \vrf/regTable[0][44] ) );
  LHQD1BWP \vrf/regTable_reg[0][45]  ( .E(n5346), .D(\vrf/N63 ), .Q(
        \vrf/regTable[0][45] ) );
  LHQD1BWP \vrf/regTable_reg[0][46]  ( .E(n5345), .D(\vrf/N64 ), .Q(
        \vrf/regTable[0][46] ) );
  LHQD1BWP \vrf/regTable_reg[0][47]  ( .E(n5345), .D(\vrf/N65 ), .Q(
        \vrf/regTable[0][47] ) );
  LHQD1BWP \vrf/regTable_reg[0][48]  ( .E(n5345), .D(\vrf/N66 ), .Q(
        \vrf/regTable[0][48] ) );
  LHQD1BWP \vrf/regTable_reg[0][49]  ( .E(n5345), .D(\vrf/N67 ), .Q(
        \vrf/regTable[0][49] ) );
  LHQD1BWP \vrf/regTable_reg[0][50]  ( .E(n5345), .D(\vrf/N68 ), .Q(
        \vrf/regTable[0][50] ) );
  LHQD1BWP \vrf/regTable_reg[0][51]  ( .E(n5345), .D(\vrf/N69 ), .Q(
        \vrf/regTable[0][51] ) );
  LHQD1BWP \vrf/regTable_reg[0][52]  ( .E(n5345), .D(\vrf/N70 ), .Q(
        \vrf/regTable[0][52] ) );
  LHQD1BWP \vrf/regTable_reg[0][53]  ( .E(n5345), .D(\vrf/N71 ), .Q(
        \vrf/regTable[0][53] ) );
  LHQD1BWP \vrf/regTable_reg[0][54]  ( .E(n5345), .D(\vrf/N72 ), .Q(
        \vrf/regTable[0][54] ) );
  LHQD1BWP \vrf/regTable_reg[0][55]  ( .E(n5345), .D(\vrf/N73 ), .Q(
        \vrf/regTable[0][55] ) );
  LHQD1BWP \vrf/regTable_reg[0][56]  ( .E(n5345), .D(\vrf/N74 ), .Q(
        \vrf/regTable[0][56] ) );
  LHQD1BWP \vrf/regTable_reg[0][57]  ( .E(n5344), .D(\vrf/N75 ), .Q(
        \vrf/regTable[0][57] ) );
  LHQD1BWP \vrf/regTable_reg[0][58]  ( .E(n5344), .D(\vrf/N76 ), .Q(
        \vrf/regTable[0][58] ) );
  LHQD1BWP \vrf/regTable_reg[0][59]  ( .E(n5344), .D(\vrf/N77 ), .Q(
        \vrf/regTable[0][59] ) );
  LHQD1BWP \vrf/regTable_reg[0][60]  ( .E(n5344), .D(\vrf/N78 ), .Q(
        \vrf/regTable[0][60] ) );
  LHQD1BWP \vrf/regTable_reg[0][61]  ( .E(n5344), .D(\vrf/N79 ), .Q(
        \vrf/regTable[0][61] ) );
  LHQD1BWP \vrf/regTable_reg[0][62]  ( .E(n5344), .D(\vrf/N80 ), .Q(
        \vrf/regTable[0][62] ) );
  LHQD1BWP \vrf/regTable_reg[0][63]  ( .E(n5344), .D(\vrf/N81 ), .Q(
        \vrf/regTable[0][63] ) );
  LHQD1BWP \vrf/regTable_reg[0][64]  ( .E(n5344), .D(\vrf/N82 ), .Q(
        \vrf/regTable[0][64] ) );
  LHQD1BWP \vrf/regTable_reg[0][65]  ( .E(n5344), .D(\vrf/N83 ), .Q(
        \vrf/regTable[0][65] ) );
  LHQD1BWP \vrf/regTable_reg[0][66]  ( .E(n5344), .D(\vrf/N84 ), .Q(
        \vrf/regTable[0][66] ) );
  LHQD1BWP \vrf/regTable_reg[0][67]  ( .E(n5344), .D(\vrf/N85 ), .Q(
        \vrf/regTable[0][67] ) );
  LHQD1BWP \vrf/regTable_reg[0][68]  ( .E(n5343), .D(\vrf/N86 ), .Q(
        \vrf/regTable[0][68] ) );
  LHQD1BWP \vrf/regTable_reg[0][69]  ( .E(n5343), .D(\vrf/N87 ), .Q(
        \vrf/regTable[0][69] ) );
  LHQD1BWP \vrf/regTable_reg[0][70]  ( .E(n5343), .D(\vrf/N88 ), .Q(
        \vrf/regTable[0][70] ) );
  LHQD1BWP \vrf/regTable_reg[0][71]  ( .E(n5343), .D(\vrf/N89 ), .Q(
        \vrf/regTable[0][71] ) );
  LHQD1BWP \vrf/regTable_reg[0][72]  ( .E(n5343), .D(\vrf/N90 ), .Q(
        \vrf/regTable[0][72] ) );
  LHQD1BWP \vrf/regTable_reg[0][73]  ( .E(n5343), .D(\vrf/N91 ), .Q(
        \vrf/regTable[0][73] ) );
  LHQD1BWP \vrf/regTable_reg[0][74]  ( .E(n5343), .D(\vrf/N92 ), .Q(
        \vrf/regTable[0][74] ) );
  LHQD1BWP \vrf/regTable_reg[0][75]  ( .E(n5343), .D(\vrf/N93 ), .Q(
        \vrf/regTable[0][75] ) );
  LHQD1BWP \vrf/regTable_reg[0][76]  ( .E(n5343), .D(\vrf/N94 ), .Q(
        \vrf/regTable[0][76] ) );
  LHQD1BWP \vrf/regTable_reg[0][77]  ( .E(n5343), .D(\vrf/N95 ), .Q(
        \vrf/regTable[0][77] ) );
  LHQD1BWP \vrf/regTable_reg[0][78]  ( .E(n5343), .D(\vrf/N96 ), .Q(
        \vrf/regTable[0][78] ) );
  LHQD1BWP \vrf/regTable_reg[0][79]  ( .E(n5342), .D(\vrf/N97 ), .Q(
        \vrf/regTable[0][79] ) );
  LHQD1BWP \vrf/regTable_reg[0][80]  ( .E(n5342), .D(\vrf/N98 ), .Q(
        \vrf/regTable[0][80] ) );
  LHQD1BWP \vrf/regTable_reg[0][81]  ( .E(n5342), .D(\vrf/N99 ), .Q(
        \vrf/regTable[0][81] ) );
  LHQD1BWP \vrf/regTable_reg[0][82]  ( .E(n5342), .D(\vrf/N100 ), .Q(
        \vrf/regTable[0][82] ) );
  LHQD1BWP \vrf/regTable_reg[0][83]  ( .E(n5342), .D(\vrf/N101 ), .Q(
        \vrf/regTable[0][83] ) );
  LHQD1BWP \vrf/regTable_reg[0][84]  ( .E(n5342), .D(\vrf/N102 ), .Q(
        \vrf/regTable[0][84] ) );
  LHQD1BWP \vrf/regTable_reg[0][85]  ( .E(n5342), .D(\vrf/N103 ), .Q(
        \vrf/regTable[0][85] ) );
  LHQD1BWP \vrf/regTable_reg[0][86]  ( .E(n5342), .D(\vrf/N104 ), .Q(
        \vrf/regTable[0][86] ) );
  LHQD1BWP \vrf/regTable_reg[0][87]  ( .E(n5342), .D(\vrf/N105 ), .Q(
        \vrf/regTable[0][87] ) );
  LHQD1BWP \vrf/regTable_reg[0][88]  ( .E(n5342), .D(\vrf/N106 ), .Q(
        \vrf/regTable[0][88] ) );
  LHQD1BWP \vrf/regTable_reg[0][89]  ( .E(n5342), .D(\vrf/N107 ), .Q(
        \vrf/regTable[0][89] ) );
  LHQD1BWP \vrf/regTable_reg[0][90]  ( .E(n5341), .D(\vrf/N108 ), .Q(
        \vrf/regTable[0][90] ) );
  LHQD1BWP \vrf/regTable_reg[0][91]  ( .E(n5341), .D(\vrf/N109 ), .Q(
        \vrf/regTable[0][91] ) );
  LHQD1BWP \vrf/regTable_reg[0][92]  ( .E(n5341), .D(\vrf/N110 ), .Q(
        \vrf/regTable[0][92] ) );
  LHQD1BWP \vrf/regTable_reg[0][93]  ( .E(n5341), .D(\vrf/N111 ), .Q(
        \vrf/regTable[0][93] ) );
  LHQD1BWP \vrf/regTable_reg[0][94]  ( .E(n5341), .D(\vrf/N112 ), .Q(
        \vrf/regTable[0][94] ) );
  LHQD1BWP \vrf/regTable_reg[0][95]  ( .E(n5341), .D(\vrf/N113 ), .Q(
        \vrf/regTable[0][95] ) );
  LHQD1BWP \vrf/regTable_reg[0][96]  ( .E(n5341), .D(\vrf/N114 ), .Q(
        \vrf/regTable[0][96] ) );
  LHQD1BWP \vrf/regTable_reg[0][97]  ( .E(n5341), .D(\vrf/N115 ), .Q(
        \vrf/regTable[0][97] ) );
  LHQD1BWP \vrf/regTable_reg[0][98]  ( .E(n5341), .D(\vrf/N116 ), .Q(
        \vrf/regTable[0][98] ) );
  LHQD1BWP \vrf/regTable_reg[0][99]  ( .E(n5341), .D(\vrf/N118 ), .Q(
        \vrf/regTable[0][99] ) );
  LHQD1BWP \vrf/regTable_reg[0][100]  ( .E(n5351), .D(\vrf/N119 ), .Q(
        \vrf/regTable[0][100] ) );
  LHQD1BWP \vrf/regTable_reg[0][101]  ( .E(n5351), .D(\vrf/N120 ), .Q(
        \vrf/regTable[0][101] ) );
  LHQD1BWP \vrf/regTable_reg[0][102]  ( .E(n5351), .D(\vrf/N121 ), .Q(
        \vrf/regTable[0][102] ) );
  LHQD1BWP \vrf/regTable_reg[0][103]  ( .E(n5351), .D(\vrf/N122 ), .Q(
        \vrf/regTable[0][103] ) );
  LHQD1BWP \vrf/regTable_reg[0][104]  ( .E(n5351), .D(\vrf/N123 ), .Q(
        \vrf/regTable[0][104] ) );
  LHQD1BWP \vrf/regTable_reg[0][105]  ( .E(n5350), .D(\vrf/N124 ), .Q(
        \vrf/regTable[0][105] ) );
  LHQD1BWP \vrf/regTable_reg[0][106]  ( .E(n5350), .D(\vrf/N125 ), .Q(
        \vrf/regTable[0][106] ) );
  LHQD1BWP \vrf/regTable_reg[0][107]  ( .E(n5350), .D(\vrf/N126 ), .Q(
        \vrf/regTable[0][107] ) );
  LHQD1BWP \vrf/regTable_reg[0][108]  ( .E(n5350), .D(\vrf/N127 ), .Q(
        \vrf/regTable[0][108] ) );
  LHQD1BWP \vrf/regTable_reg[0][109]  ( .E(n5350), .D(\vrf/N128 ), .Q(
        \vrf/regTable[0][109] ) );
  LHQD1BWP \vrf/regTable_reg[0][110]  ( .E(n5350), .D(\vrf/N129 ), .Q(
        \vrf/regTable[0][110] ) );
  LHQD1BWP \vrf/regTable_reg[0][111]  ( .E(n5350), .D(\vrf/N130 ), .Q(
        \vrf/regTable[0][111] ) );
  LHQD1BWP \vrf/regTable_reg[0][112]  ( .E(n5350), .D(\vrf/N131 ), .Q(
        \vrf/regTable[0][112] ) );
  LHQD1BWP \vrf/regTable_reg[0][113]  ( .E(n5350), .D(\vrf/N132 ), .Q(
        \vrf/regTable[0][113] ) );
  LHQD1BWP \vrf/regTable_reg[0][114]  ( .E(n5350), .D(\vrf/N133 ), .Q(
        \vrf/regTable[0][114] ) );
  LHQD1BWP \vrf/regTable_reg[0][115]  ( .E(n5350), .D(\vrf/N134 ), .Q(
        \vrf/regTable[0][115] ) );
  LHQD1BWP \vrf/regTable_reg[0][116]  ( .E(n5349), .D(\vrf/N135 ), .Q(
        \vrf/regTable[0][116] ) );
  LHQD1BWP \vrf/regTable_reg[0][117]  ( .E(n5349), .D(\vrf/N136 ), .Q(
        \vrf/regTable[0][117] ) );
  LHQD1BWP \vrf/regTable_reg[0][118]  ( .E(n5349), .D(\vrf/N137 ), .Q(
        \vrf/regTable[0][118] ) );
  LHQD1BWP \vrf/regTable_reg[0][119]  ( .E(n5349), .D(\vrf/N138 ), .Q(
        \vrf/regTable[0][119] ) );
  LHQD1BWP \vrf/regTable_reg[0][120]  ( .E(n5349), .D(\vrf/N139 ), .Q(
        \vrf/regTable[0][120] ) );
  LHQD1BWP \vrf/regTable_reg[0][121]  ( .E(n5349), .D(\vrf/N140 ), .Q(
        \vrf/regTable[0][121] ) );
  LHQD1BWP \vrf/regTable_reg[0][122]  ( .E(n5349), .D(\vrf/N141 ), .Q(
        \vrf/regTable[0][122] ) );
  LHQD1BWP \vrf/regTable_reg[0][123]  ( .E(n5349), .D(\vrf/N142 ), .Q(
        \vrf/regTable[0][123] ) );
  LHQD1BWP \vrf/regTable_reg[0][124]  ( .E(n5349), .D(\vrf/N143 ), .Q(
        \vrf/regTable[0][124] ) );
  LHQD1BWP \vrf/regTable_reg[0][125]  ( .E(n5349), .D(\vrf/N144 ), .Q(
        \vrf/regTable[0][125] ) );
  LHQD1BWP \vrf/regTable_reg[0][126]  ( .E(n5349), .D(\vrf/N145 ), .Q(
        \vrf/regTable[0][126] ) );
  LHQD1BWP \vrf/regTable_reg[0][127]  ( .E(n5348), .D(\vrf/N146 ), .Q(
        \vrf/regTable[0][127] ) );
  LHQD1BWP \vrf/regTable_reg[0][128]  ( .E(n5351), .D(\vrf/N147 ), .Q(
        \vrf/regTable[0][128] ) );
  LHQD1BWP \vrf/regTable_reg[0][129]  ( .E(n5351), .D(\vrf/N148 ), .Q(
        \vrf/regTable[0][129] ) );
  LHQD1BWP \vrf/regTable_reg[0][130]  ( .E(n5351), .D(\vrf/N149 ), .Q(
        \vrf/regTable[0][130] ) );
  LHQD1BWP \vrf/regTable_reg[0][131]  ( .E(n5351), .D(\vrf/N150 ), .Q(
        \vrf/regTable[0][131] ) );
  LHQD1BWP \vrf/regTable_reg[0][132]  ( .E(n5351), .D(\vrf/N151 ), .Q(
        \vrf/regTable[0][132] ) );
  LHQD1BWP \vrf/regTable_reg[0][133]  ( .E(n5351), .D(\vrf/N152 ), .Q(
        \vrf/regTable[0][133] ) );
  LHQD1BWP \vrf/regTable_reg[0][134]  ( .E(n5352), .D(\vrf/N153 ), .Q(
        \vrf/regTable[0][134] ) );
  LHQD1BWP \vrf/regTable_reg[0][135]  ( .E(n5352), .D(\vrf/N154 ), .Q(
        \vrf/regTable[0][135] ) );
  LHQD1BWP \vrf/regTable_reg[0][136]  ( .E(n5352), .D(\vrf/N155 ), .Q(
        \vrf/regTable[0][136] ) );
  LHQD1BWP \vrf/regTable_reg[0][137]  ( .E(n5352), .D(\vrf/N156 ), .Q(
        \vrf/regTable[0][137] ) );
  LHQD1BWP \vrf/regTable_reg[0][138]  ( .E(n5352), .D(\vrf/N157 ), .Q(
        \vrf/regTable[0][138] ) );
  LHQD1BWP \vrf/regTable_reg[0][139]  ( .E(n5352), .D(\vrf/N158 ), .Q(
        \vrf/regTable[0][139] ) );
  LHQD1BWP \vrf/regTable_reg[0][140]  ( .E(n5352), .D(\vrf/N159 ), .Q(
        \vrf/regTable[0][140] ) );
  LHQD1BWP \vrf/regTable_reg[0][141]  ( .E(n5352), .D(\vrf/N160 ), .Q(
        \vrf/regTable[0][141] ) );
  LHQD1BWP \vrf/regTable_reg[0][142]  ( .E(n5352), .D(\vrf/N161 ), .Q(
        \vrf/regTable[0][142] ) );
  LHQD1BWP \vrf/regTable_reg[0][143]  ( .E(n5352), .D(\vrf/N162 ), .Q(
        \vrf/regTable[0][143] ) );
  LHQD1BWP \vrf/regTable_reg[0][144]  ( .E(n5352), .D(\vrf/N163 ), .Q(
        \vrf/regTable[0][144] ) );
  LHQD1BWP \vrf/regTable_reg[0][145]  ( .E(n5352), .D(\vrf/N164 ), .Q(
        \vrf/regTable[0][145] ) );
  LHQD1BWP \vrf/regTable_reg[0][146]  ( .E(n5353), .D(\vrf/N165 ), .Q(
        \vrf/regTable[0][146] ) );
  LHQD1BWP \vrf/regTable_reg[0][147]  ( .E(n5353), .D(\vrf/N166 ), .Q(
        \vrf/regTable[0][147] ) );
  LHQD1BWP \vrf/regTable_reg[0][148]  ( .E(n5353), .D(\vrf/N167 ), .Q(
        \vrf/regTable[0][148] ) );
  LHQD1BWP \vrf/regTable_reg[0][149]  ( .E(n5353), .D(\vrf/N168 ), .Q(
        \vrf/regTable[0][149] ) );
  LHQD1BWP \vrf/regTable_reg[0][150]  ( .E(n5353), .D(\vrf/N169 ), .Q(
        \vrf/regTable[0][150] ) );
  LHQD1BWP \vrf/regTable_reg[0][151]  ( .E(n5353), .D(\vrf/N170 ), .Q(
        \vrf/regTable[0][151] ) );
  LHQD1BWP \vrf/regTable_reg[0][152]  ( .E(n5353), .D(\vrf/N171 ), .Q(
        \vrf/regTable[0][152] ) );
  LHQD1BWP \vrf/regTable_reg[0][153]  ( .E(n5353), .D(\vrf/N172 ), .Q(
        \vrf/regTable[0][153] ) );
  LHQD1BWP \vrf/regTable_reg[0][154]  ( .E(n5353), .D(\vrf/N173 ), .Q(
        \vrf/regTable[0][154] ) );
  LHQD1BWP \vrf/regTable_reg[0][155]  ( .E(n5353), .D(\vrf/N174 ), .Q(
        \vrf/regTable[0][155] ) );
  LHQD1BWP \vrf/regTable_reg[0][156]  ( .E(n5353), .D(\vrf/N175 ), .Q(
        \vrf/regTable[0][156] ) );
  LHQD1BWP \vrf/regTable_reg[0][157]  ( .E(n5353), .D(\vrf/N176 ), .Q(
        \vrf/regTable[0][157] ) );
  LHQD1BWP \vrf/regTable_reg[0][158]  ( .E(n5354), .D(\vrf/N177 ), .Q(
        \vrf/regTable[0][158] ) );
  LHQD1BWP \vrf/regTable_reg[0][159]  ( .E(n5354), .D(\vrf/N178 ), .Q(
        \vrf/regTable[0][159] ) );
  LHQD1BWP \vrf/regTable_reg[0][160]  ( .E(n5354), .D(\vrf/N179 ), .Q(
        \vrf/regTable[0][160] ) );
  LHQD1BWP \vrf/regTable_reg[0][161]  ( .E(n5354), .D(\vrf/N180 ), .Q(
        \vrf/regTable[0][161] ) );
  LHQD1BWP \vrf/regTable_reg[0][162]  ( .E(n5354), .D(\vrf/N181 ), .Q(
        \vrf/regTable[0][162] ) );
  LHQD1BWP \vrf/regTable_reg[0][163]  ( .E(n5354), .D(\vrf/N182 ), .Q(
        \vrf/regTable[0][163] ) );
  LHQD1BWP \vrf/regTable_reg[0][164]  ( .E(n5354), .D(\vrf/N183 ), .Q(
        \vrf/regTable[0][164] ) );
  LHQD1BWP \vrf/regTable_reg[0][165]  ( .E(n5354), .D(\vrf/N184 ), .Q(
        \vrf/regTable[0][165] ) );
  LHQD1BWP \vrf/regTable_reg[0][166]  ( .E(n5354), .D(\vrf/N185 ), .Q(
        \vrf/regTable[0][166] ) );
  LHQD1BWP \vrf/regTable_reg[0][167]  ( .E(n5354), .D(\vrf/N186 ), .Q(
        \vrf/regTable[0][167] ) );
  LHQD1BWP \vrf/regTable_reg[0][168]  ( .E(n5354), .D(\vrf/N187 ), .Q(
        \vrf/regTable[0][168] ) );
  LHQD1BWP \vrf/regTable_reg[0][169]  ( .E(n5354), .D(\vrf/N188 ), .Q(
        \vrf/regTable[0][169] ) );
  LHQD1BWP \vrf/regTable_reg[0][170]  ( .E(n5355), .D(\vrf/N189 ), .Q(
        \vrf/regTable[0][170] ) );
  LHQD1BWP \vrf/regTable_reg[0][171]  ( .E(n5355), .D(\vrf/N190 ), .Q(
        \vrf/regTable[0][171] ) );
  LHQD1BWP \vrf/regTable_reg[0][172]  ( .E(n5355), .D(\vrf/N191 ), .Q(
        \vrf/regTable[0][172] ) );
  LHQD1BWP \vrf/regTable_reg[0][173]  ( .E(n5355), .D(\vrf/N192 ), .Q(
        \vrf/regTable[0][173] ) );
  LHQD1BWP \vrf/regTable_reg[0][174]  ( .E(n5355), .D(\vrf/N193 ), .Q(
        \vrf/regTable[0][174] ) );
  LHQD1BWP \vrf/regTable_reg[0][175]  ( .E(n5355), .D(\vrf/N194 ), .Q(
        \vrf/regTable[0][175] ) );
  LHQD1BWP \vrf/regTable_reg[0][176]  ( .E(n5355), .D(\vrf/N195 ), .Q(
        \vrf/regTable[0][176] ) );
  LHQD1BWP \vrf/regTable_reg[0][177]  ( .E(n5355), .D(\vrf/N196 ), .Q(
        \vrf/regTable[0][177] ) );
  LHQD1BWP \vrf/regTable_reg[0][178]  ( .E(n5355), .D(\vrf/N197 ), .Q(
        \vrf/regTable[0][178] ) );
  LHQD1BWP \vrf/regTable_reg[0][179]  ( .E(n5355), .D(\vrf/N198 ), .Q(
        \vrf/regTable[0][179] ) );
  LHQD1BWP \vrf/regTable_reg[0][180]  ( .E(n5355), .D(\vrf/N199 ), .Q(
        \vrf/regTable[0][180] ) );
  LHQD1BWP \vrf/regTable_reg[0][181]  ( .E(n5355), .D(\vrf/N200 ), .Q(
        \vrf/regTable[0][181] ) );
  LHQD1BWP \vrf/regTable_reg[0][182]  ( .E(n5356), .D(\vrf/N201 ), .Q(
        \vrf/regTable[0][182] ) );
  LHQD1BWP \vrf/regTable_reg[0][183]  ( .E(n5356), .D(\vrf/N202 ), .Q(
        \vrf/regTable[0][183] ) );
  LHQD1BWP \vrf/regTable_reg[0][184]  ( .E(n5356), .D(\vrf/N203 ), .Q(
        \vrf/regTable[0][184] ) );
  LHQD1BWP \vrf/regTable_reg[0][185]  ( .E(n5356), .D(\vrf/N204 ), .Q(
        \vrf/regTable[0][185] ) );
  LHQD1BWP \vrf/regTable_reg[0][186]  ( .E(n5356), .D(\vrf/N205 ), .Q(
        \vrf/regTable[0][186] ) );
  LHQD1BWP \vrf/regTable_reg[0][187]  ( .E(n5356), .D(\vrf/N206 ), .Q(
        \vrf/regTable[0][187] ) );
  LHQD1BWP \vrf/regTable_reg[0][188]  ( .E(n5356), .D(\vrf/N207 ), .Q(
        \vrf/regTable[0][188] ) );
  LHQD1BWP \vrf/regTable_reg[0][189]  ( .E(n5356), .D(\vrf/N208 ), .Q(
        \vrf/regTable[0][189] ) );
  LHQD1BWP \vrf/regTable_reg[0][190]  ( .E(n5356), .D(\vrf/N209 ), .Q(
        \vrf/regTable[0][190] ) );
  LHQD1BWP \vrf/regTable_reg[0][191]  ( .E(n5356), .D(\vrf/N210 ), .Q(
        \vrf/regTable[0][191] ) );
  LHQD1BWP \vrf/regTable_reg[0][192]  ( .E(n5356), .D(\vrf/N211 ), .Q(
        \vrf/regTable[0][192] ) );
  LHQD1BWP \vrf/regTable_reg[0][193]  ( .E(n5356), .D(\vrf/N212 ), .Q(
        \vrf/regTable[0][193] ) );
  LHQD1BWP \vrf/regTable_reg[0][194]  ( .E(n5357), .D(\vrf/N213 ), .Q(
        \vrf/regTable[0][194] ) );
  LHQD1BWP \vrf/regTable_reg[0][195]  ( .E(n5357), .D(\vrf/N214 ), .Q(
        \vrf/regTable[0][195] ) );
  LHQD1BWP \vrf/regTable_reg[0][196]  ( .E(n5357), .D(\vrf/N215 ), .Q(
        \vrf/regTable[0][196] ) );
  LHQD1BWP \vrf/regTable_reg[0][197]  ( .E(n5357), .D(\vrf/N216 ), .Q(
        \vrf/regTable[0][197] ) );
  LHQD1BWP \vrf/regTable_reg[0][198]  ( .E(n5357), .D(\vrf/N218 ), .Q(
        \vrf/regTable[0][198] ) );
  LHQD1BWP \vrf/regTable_reg[0][199]  ( .E(n5357), .D(\vrf/N219 ), .Q(
        \vrf/regTable[0][199] ) );
  LHQD1BWP \vrf/regTable_reg[0][200]  ( .E(n5357), .D(\vrf/N220 ), .Q(
        \vrf/regTable[0][200] ) );
  LHQD1BWP \vrf/regTable_reg[0][201]  ( .E(n5357), .D(\vrf/N221 ), .Q(
        \vrf/regTable[0][201] ) );
  LHQD1BWP \vrf/regTable_reg[0][202]  ( .E(n5357), .D(\vrf/N222 ), .Q(
        \vrf/regTable[0][202] ) );
  LHQD1BWP \vrf/regTable_reg[0][203]  ( .E(n5357), .D(\vrf/N223 ), .Q(
        \vrf/regTable[0][203] ) );
  LHQD1BWP \vrf/regTable_reg[0][204]  ( .E(n5357), .D(\vrf/N224 ), .Q(
        \vrf/regTable[0][204] ) );
  LHQD1BWP \vrf/regTable_reg[0][205]  ( .E(n5357), .D(\vrf/N225 ), .Q(
        \vrf/regTable[0][205] ) );
  LHQD1BWP \vrf/regTable_reg[0][206]  ( .E(n5358), .D(\vrf/N226 ), .Q(
        \vrf/regTable[0][206] ) );
  LHQD1BWP \vrf/regTable_reg[0][207]  ( .E(n5358), .D(\vrf/N227 ), .Q(
        \vrf/regTable[0][207] ) );
  LHQD1BWP \vrf/regTable_reg[0][208]  ( .E(n5358), .D(\vrf/N228 ), .Q(
        \vrf/regTable[0][208] ) );
  LHQD1BWP \vrf/regTable_reg[0][209]  ( .E(n5358), .D(\vrf/N229 ), .Q(
        \vrf/regTable[0][209] ) );
  LHQD1BWP \vrf/regTable_reg[0][210]  ( .E(n5358), .D(\vrf/N230 ), .Q(
        \vrf/regTable[0][210] ) );
  LHQD1BWP \vrf/regTable_reg[0][211]  ( .E(n5358), .D(\vrf/N231 ), .Q(
        \vrf/regTable[0][211] ) );
  LHQD1BWP \vrf/regTable_reg[0][212]  ( .E(n5358), .D(\vrf/N232 ), .Q(
        \vrf/regTable[0][212] ) );
  LHQD1BWP \vrf/regTable_reg[0][213]  ( .E(n5358), .D(\vrf/N233 ), .Q(
        \vrf/regTable[0][213] ) );
  LHQD1BWP \vrf/regTable_reg[0][214]  ( .E(n5358), .D(\vrf/N234 ), .Q(
        \vrf/regTable[0][214] ) );
  LHQD1BWP \vrf/regTable_reg[0][215]  ( .E(n5358), .D(\vrf/N235 ), .Q(
        \vrf/regTable[0][215] ) );
  LHQD1BWP \vrf/regTable_reg[0][216]  ( .E(n5358), .D(\vrf/N236 ), .Q(
        \vrf/regTable[0][216] ) );
  LHQD1BWP \vrf/regTable_reg[0][217]  ( .E(n5358), .D(\vrf/N237 ), .Q(
        \vrf/regTable[0][217] ) );
  LHQD1BWP \vrf/regTable_reg[0][218]  ( .E(n5359), .D(\vrf/N238 ), .Q(
        \vrf/regTable[0][218] ) );
  LHQD1BWP \vrf/regTable_reg[0][219]  ( .E(n5359), .D(\vrf/N239 ), .Q(
        \vrf/regTable[0][219] ) );
  LHQD1BWP \vrf/regTable_reg[0][220]  ( .E(n5359), .D(\vrf/N240 ), .Q(
        \vrf/regTable[0][220] ) );
  LHQD1BWP \vrf/regTable_reg[0][221]  ( .E(n5359), .D(\vrf/N241 ), .Q(
        \vrf/regTable[0][221] ) );
  LHQD1BWP \vrf/regTable_reg[0][222]  ( .E(n5359), .D(\vrf/N242 ), .Q(
        \vrf/regTable[0][222] ) );
  LHQD1BWP \vrf/regTable_reg[0][223]  ( .E(n5359), .D(\vrf/N243 ), .Q(
        \vrf/regTable[0][223] ) );
  LHQD1BWP \vrf/regTable_reg[0][224]  ( .E(n5359), .D(\vrf/N244 ), .Q(
        \vrf/regTable[0][224] ) );
  LHQD1BWP \vrf/regTable_reg[0][225]  ( .E(n5359), .D(\vrf/N245 ), .Q(
        \vrf/regTable[0][225] ) );
  LHQD1BWP \vrf/regTable_reg[0][226]  ( .E(n5359), .D(\vrf/N246 ), .Q(
        \vrf/regTable[0][226] ) );
  LHQD1BWP \vrf/regTable_reg[0][227]  ( .E(n5359), .D(\vrf/N247 ), .Q(
        \vrf/regTable[0][227] ) );
  LHQD1BWP \vrf/regTable_reg[0][228]  ( .E(n5359), .D(\vrf/N248 ), .Q(
        \vrf/regTable[0][228] ) );
  LHQD1BWP \vrf/regTable_reg[0][229]  ( .E(n5359), .D(\vrf/N249 ), .Q(
        \vrf/regTable[0][229] ) );
  LHQD1BWP \vrf/regTable_reg[0][230]  ( .E(n5360), .D(\vrf/N250 ), .Q(
        \vrf/regTable[0][230] ) );
  LHQD1BWP \vrf/regTable_reg[0][231]  ( .E(n5360), .D(\vrf/N251 ), .Q(
        \vrf/regTable[0][231] ) );
  LHQD1BWP \vrf/regTable_reg[0][232]  ( .E(n5360), .D(\vrf/N252 ), .Q(
        \vrf/regTable[0][232] ) );
  LHQD1BWP \vrf/regTable_reg[0][233]  ( .E(n5360), .D(\vrf/N253 ), .Q(
        \vrf/regTable[0][233] ) );
  LHQD1BWP \vrf/regTable_reg[0][234]  ( .E(n5360), .D(\vrf/N254 ), .Q(
        \vrf/regTable[0][234] ) );
  LHQD1BWP \vrf/regTable_reg[0][235]  ( .E(n5360), .D(\vrf/N255 ), .Q(
        \vrf/regTable[0][235] ) );
  LHQD1BWP \vrf/regTable_reg[0][236]  ( .E(n5360), .D(\vrf/N256 ), .Q(
        \vrf/regTable[0][236] ) );
  LHQD1BWP \vrf/regTable_reg[0][237]  ( .E(n5360), .D(\vrf/N257 ), .Q(
        \vrf/regTable[0][237] ) );
  LHQD1BWP \vrf/regTable_reg[0][238]  ( .E(n5360), .D(\vrf/N258 ), .Q(
        \vrf/regTable[0][238] ) );
  LHQD1BWP \vrf/regTable_reg[0][239]  ( .E(n5360), .D(\vrf/N259 ), .Q(
        \vrf/regTable[0][239] ) );
  LHQD1BWP \vrf/regTable_reg[0][240]  ( .E(n5360), .D(\vrf/N260 ), .Q(
        \vrf/regTable[0][240] ) );
  LHQD1BWP \vrf/regTable_reg[0][241]  ( .E(n5360), .D(\vrf/N261 ), .Q(
        \vrf/regTable[0][241] ) );
  LHQD1BWP \vrf/regTable_reg[0][242]  ( .E(n5361), .D(\vrf/N262 ), .Q(
        \vrf/regTable[0][242] ) );
  LHQD1BWP \vrf/regTable_reg[0][243]  ( .E(n5361), .D(\vrf/N263 ), .Q(
        \vrf/regTable[0][243] ) );
  LHQD1BWP \vrf/regTable_reg[0][244]  ( .E(n5361), .D(\vrf/N264 ), .Q(
        \vrf/regTable[0][244] ) );
  LHQD1BWP \vrf/regTable_reg[0][245]  ( .E(n5361), .D(\vrf/N265 ), .Q(
        \vrf/regTable[0][245] ) );
  LHQD1BWP \vrf/regTable_reg[0][246]  ( .E(n5361), .D(\vrf/N266 ), .Q(
        \vrf/regTable[0][246] ) );
  LHQD1BWP \vrf/regTable_reg[0][247]  ( .E(n5361), .D(\vrf/N267 ), .Q(
        \vrf/regTable[0][247] ) );
  LHQD1BWP \vrf/regTable_reg[0][248]  ( .E(n5361), .D(\vrf/N268 ), .Q(
        \vrf/regTable[0][248] ) );
  LHQD1BWP \vrf/regTable_reg[0][249]  ( .E(n5361), .D(\vrf/N269 ), .Q(
        \vrf/regTable[0][249] ) );
  LHQD1BWP \vrf/regTable_reg[0][250]  ( .E(n5361), .D(\vrf/N270 ), .Q(
        \vrf/regTable[0][250] ) );
  LHQD1BWP \vrf/regTable_reg[0][251]  ( .E(n5361), .D(\vrf/N271 ), .Q(
        \vrf/regTable[0][251] ) );
  LHQD1BWP \vrf/regTable_reg[0][252]  ( .E(n5361), .D(\vrf/N272 ), .Q(
        \vrf/regTable[0][252] ) );
  LHQD1BWP \vrf/regTable_reg[0][253]  ( .E(n5361), .D(\vrf/N273 ), .Q(
        \vrf/regTable[0][253] ) );
  LHQD1BWP \vrf/regTable_reg[7][15]  ( .E(n5124), .D(\vrf/N33 ), .Q(
        \vrf/regTable[7][15] ) );
  LHQD1BWP \vrf/regTable_reg[7][16]  ( .E(n5124), .D(\vrf/N34 ), .Q(
        \vrf/regTable[7][16] ) );
  LHQD1BWP \vrf/regTable_reg[7][254]  ( .E(n5124), .D(\vrf/N274 ), .Q(
        \vrf/regTable[7][254] ) );
  LHQD1BWP \vrf/regTable_reg[7][255]  ( .E(n5124), .D(\vrf/N275 ), .Q(
        \vrf/regTable[7][255] ) );
  LHQD1BWP \vrf/regTable_reg[3][15]  ( .E(n5260), .D(\vrf/N33 ), .Q(
        \vrf/regTable[3][15] ) );
  LHQD1BWP \vrf/regTable_reg[3][16]  ( .E(n5260), .D(\vrf/N34 ), .Q(
        \vrf/regTable[3][16] ) );
  LHQD1BWP \vrf/regTable_reg[3][254]  ( .E(n5260), .D(\vrf/N274 ), .Q(
        \vrf/regTable[3][254] ) );
  LHQD1BWP \vrf/regTable_reg[3][255]  ( .E(n5260), .D(\vrf/N275 ), .Q(
        \vrf/regTable[3][255] ) );
  LHQD1BWP \vrf/regTable_reg[7][0]  ( .E(n5113), .D(\vrf/N18 ), .Q(
        \vrf/regTable[7][0] ) );
  LHQD1BWP \vrf/regTable_reg[7][1]  ( .E(n5110), .D(\vrf/N19 ), .Q(
        \vrf/regTable[7][1] ) );
  LHQD1BWP \vrf/regTable_reg[7][2]  ( .E(n5109), .D(\vrf/N20 ), .Q(
        \vrf/regTable[7][2] ) );
  LHQD1BWP \vrf/regTable_reg[7][3]  ( .E(n5108), .D(\vrf/N21 ), .Q(
        \vrf/regTable[7][3] ) );
  LHQD1BWP \vrf/regTable_reg[7][4]  ( .E(n5107), .D(\vrf/N22 ), .Q(
        \vrf/regTable[7][4] ) );
  LHQD1BWP \vrf/regTable_reg[7][5]  ( .E(n5106), .D(\vrf/N23 ), .Q(
        \vrf/regTable[7][5] ) );
  LHQD1BWP \vrf/regTable_reg[7][6]  ( .E(n5105), .D(\vrf/N24 ), .Q(
        \vrf/regTable[7][6] ) );
  LHQD1BWP \vrf/regTable_reg[7][7]  ( .E(n5104), .D(\vrf/N25 ), .Q(
        \vrf/regTable[7][7] ) );
  LHQD1BWP \vrf/regTable_reg[7][8]  ( .E(n5103), .D(\vrf/N26 ), .Q(
        \vrf/regTable[7][8] ) );
  LHQD1BWP \vrf/regTable_reg[7][9]  ( .E(n5103), .D(\vrf/N27 ), .Q(
        \vrf/regTable[7][9] ) );
  LHQD1BWP \vrf/regTable_reg[7][10]  ( .E(n5112), .D(\vrf/N28 ), .Q(
        \vrf/regTable[7][10] ) );
  LHQD1BWP \vrf/regTable_reg[7][11]  ( .E(n5111), .D(\vrf/N29 ), .Q(
        \vrf/regTable[7][11] ) );
  LHQD1BWP \vrf/regTable_reg[7][12]  ( .E(n5110), .D(\vrf/N30 ), .Q(
        \vrf/regTable[7][12] ) );
  LHQD1BWP \vrf/regTable_reg[7][13]  ( .E(n5110), .D(\vrf/N31 ), .Q(
        \vrf/regTable[7][13] ) );
  LHQD1BWP \vrf/regTable_reg[7][14]  ( .E(n5110), .D(\vrf/N32 ), .Q(
        \vrf/regTable[7][14] ) );
  LHQD1BWP \vrf/regTable_reg[7][17]  ( .E(n5110), .D(\vrf/N35 ), .Q(
        \vrf/regTable[7][17] ) );
  LHQD1BWP \vrf/regTable_reg[7][18]  ( .E(n5110), .D(\vrf/N36 ), .Q(
        \vrf/regTable[7][18] ) );
  LHQD1BWP \vrf/regTable_reg[7][19]  ( .E(n5110), .D(\vrf/N37 ), .Q(
        \vrf/regTable[7][19] ) );
  LHQD1BWP \vrf/regTable_reg[7][20]  ( .E(n5110), .D(\vrf/N38 ), .Q(
        \vrf/regTable[7][20] ) );
  LHQD1BWP \vrf/regTable_reg[7][21]  ( .E(n5110), .D(\vrf/N39 ), .Q(
        \vrf/regTable[7][21] ) );
  LHQD1BWP \vrf/regTable_reg[7][22]  ( .E(n5110), .D(\vrf/N40 ), .Q(
        \vrf/regTable[7][22] ) );
  LHQD1BWP \vrf/regTable_reg[7][23]  ( .E(n5110), .D(\vrf/N41 ), .Q(
        \vrf/regTable[7][23] ) );
  LHQD1BWP \vrf/regTable_reg[7][24]  ( .E(n5109), .D(\vrf/N42 ), .Q(
        \vrf/regTable[7][24] ) );
  LHQD1BWP \vrf/regTable_reg[7][25]  ( .E(n5109), .D(\vrf/N43 ), .Q(
        \vrf/regTable[7][25] ) );
  LHQD1BWP \vrf/regTable_reg[7][26]  ( .E(n5109), .D(\vrf/N44 ), .Q(
        \vrf/regTable[7][26] ) );
  LHQD1BWP \vrf/regTable_reg[7][27]  ( .E(n5109), .D(\vrf/N45 ), .Q(
        \vrf/regTable[7][27] ) );
  LHQD1BWP \vrf/regTable_reg[7][28]  ( .E(n5109), .D(\vrf/N46 ), .Q(
        \vrf/regTable[7][28] ) );
  LHQD1BWP \vrf/regTable_reg[7][29]  ( .E(n5109), .D(\vrf/N47 ), .Q(
        \vrf/regTable[7][29] ) );
  LHQD1BWP \vrf/regTable_reg[7][30]  ( .E(n5109), .D(\vrf/N48 ), .Q(
        \vrf/regTable[7][30] ) );
  LHQD1BWP \vrf/regTable_reg[7][31]  ( .E(n5109), .D(\vrf/N49 ), .Q(
        \vrf/regTable[7][31] ) );
  LHQD1BWP \vrf/regTable_reg[7][32]  ( .E(n5109), .D(\vrf/N50 ), .Q(
        \vrf/regTable[7][32] ) );
  LHQD1BWP \vrf/regTable_reg[7][33]  ( .E(n5109), .D(\vrf/N51 ), .Q(
        \vrf/regTable[7][33] ) );
  LHQD1BWP \vrf/regTable_reg[7][34]  ( .E(n5109), .D(\vrf/N52 ), .Q(
        \vrf/regTable[7][34] ) );
  LHQD1BWP \vrf/regTable_reg[7][35]  ( .E(n5108), .D(\vrf/N53 ), .Q(
        \vrf/regTable[7][35] ) );
  LHQD1BWP \vrf/regTable_reg[7][36]  ( .E(n5108), .D(\vrf/N54 ), .Q(
        \vrf/regTable[7][36] ) );
  LHQD1BWP \vrf/regTable_reg[7][37]  ( .E(n5108), .D(\vrf/N55 ), .Q(
        \vrf/regTable[7][37] ) );
  LHQD1BWP \vrf/regTable_reg[7][38]  ( .E(n5108), .D(\vrf/N56 ), .Q(
        \vrf/regTable[7][38] ) );
  LHQD1BWP \vrf/regTable_reg[7][39]  ( .E(n5108), .D(\vrf/N57 ), .Q(
        \vrf/regTable[7][39] ) );
  LHQD1BWP \vrf/regTable_reg[7][40]  ( .E(n5108), .D(\vrf/N58 ), .Q(
        \vrf/regTable[7][40] ) );
  LHQD1BWP \vrf/regTable_reg[7][41]  ( .E(n5108), .D(\vrf/N59 ), .Q(
        \vrf/regTable[7][41] ) );
  LHQD1BWP \vrf/regTable_reg[7][42]  ( .E(n5108), .D(\vrf/N60 ), .Q(
        \vrf/regTable[7][42] ) );
  LHQD1BWP \vrf/regTable_reg[7][43]  ( .E(n5108), .D(\vrf/N61 ), .Q(
        \vrf/regTable[7][43] ) );
  LHQD1BWP \vrf/regTable_reg[7][44]  ( .E(n5108), .D(\vrf/N62 ), .Q(
        \vrf/regTable[7][44] ) );
  LHQD1BWP \vrf/regTable_reg[7][45]  ( .E(n5108), .D(\vrf/N63 ), .Q(
        \vrf/regTable[7][45] ) );
  LHQD1BWP \vrf/regTable_reg[7][46]  ( .E(n5107), .D(\vrf/N64 ), .Q(
        \vrf/regTable[7][46] ) );
  LHQD1BWP \vrf/regTable_reg[7][47]  ( .E(n5107), .D(\vrf/N65 ), .Q(
        \vrf/regTable[7][47] ) );
  LHQD1BWP \vrf/regTable_reg[7][48]  ( .E(n5107), .D(\vrf/N66 ), .Q(
        \vrf/regTable[7][48] ) );
  LHQD1BWP \vrf/regTable_reg[7][49]  ( .E(n5107), .D(\vrf/N67 ), .Q(
        \vrf/regTable[7][49] ) );
  LHQD1BWP \vrf/regTable_reg[7][50]  ( .E(n5107), .D(\vrf/N68 ), .Q(
        \vrf/regTable[7][50] ) );
  LHQD1BWP \vrf/regTable_reg[7][51]  ( .E(n5107), .D(\vrf/N69 ), .Q(
        \vrf/regTable[7][51] ) );
  LHQD1BWP \vrf/regTable_reg[7][52]  ( .E(n5107), .D(\vrf/N70 ), .Q(
        \vrf/regTable[7][52] ) );
  LHQD1BWP \vrf/regTable_reg[7][53]  ( .E(n5107), .D(\vrf/N71 ), .Q(
        \vrf/regTable[7][53] ) );
  LHQD1BWP \vrf/regTable_reg[7][54]  ( .E(n5107), .D(\vrf/N72 ), .Q(
        \vrf/regTable[7][54] ) );
  LHQD1BWP \vrf/regTable_reg[7][55]  ( .E(n5107), .D(\vrf/N73 ), .Q(
        \vrf/regTable[7][55] ) );
  LHQD1BWP \vrf/regTable_reg[7][56]  ( .E(n5107), .D(\vrf/N74 ), .Q(
        \vrf/regTable[7][56] ) );
  LHQD1BWP \vrf/regTable_reg[7][57]  ( .E(n5106), .D(\vrf/N75 ), .Q(
        \vrf/regTable[7][57] ) );
  LHQD1BWP \vrf/regTable_reg[7][58]  ( .E(n5106), .D(\vrf/N76 ), .Q(
        \vrf/regTable[7][58] ) );
  LHQD1BWP \vrf/regTable_reg[7][59]  ( .E(n5106), .D(\vrf/N77 ), .Q(
        \vrf/regTable[7][59] ) );
  LHQD1BWP \vrf/regTable_reg[7][60]  ( .E(n5106), .D(\vrf/N78 ), .Q(
        \vrf/regTable[7][60] ) );
  LHQD1BWP \vrf/regTable_reg[7][61]  ( .E(n5106), .D(\vrf/N79 ), .Q(
        \vrf/regTable[7][61] ) );
  LHQD1BWP \vrf/regTable_reg[7][62]  ( .E(n5106), .D(\vrf/N80 ), .Q(
        \vrf/regTable[7][62] ) );
  LHQD1BWP \vrf/regTable_reg[7][63]  ( .E(n5106), .D(\vrf/N81 ), .Q(
        \vrf/regTable[7][63] ) );
  LHQD1BWP \vrf/regTable_reg[7][64]  ( .E(n5106), .D(\vrf/N82 ), .Q(
        \vrf/regTable[7][64] ) );
  LHQD1BWP \vrf/regTable_reg[7][65]  ( .E(n5106), .D(\vrf/N83 ), .Q(
        \vrf/regTable[7][65] ) );
  LHQD1BWP \vrf/regTable_reg[7][66]  ( .E(n5106), .D(\vrf/N84 ), .Q(
        \vrf/regTable[7][66] ) );
  LHQD1BWP \vrf/regTable_reg[7][67]  ( .E(n5106), .D(\vrf/N85 ), .Q(
        \vrf/regTable[7][67] ) );
  LHQD1BWP \vrf/regTable_reg[7][68]  ( .E(n5105), .D(\vrf/N86 ), .Q(
        \vrf/regTable[7][68] ) );
  LHQD1BWP \vrf/regTable_reg[7][69]  ( .E(n5105), .D(\vrf/N87 ), .Q(
        \vrf/regTable[7][69] ) );
  LHQD1BWP \vrf/regTable_reg[7][70]  ( .E(n5105), .D(\vrf/N88 ), .Q(
        \vrf/regTable[7][70] ) );
  LHQD1BWP \vrf/regTable_reg[7][71]  ( .E(n5105), .D(\vrf/N89 ), .Q(
        \vrf/regTable[7][71] ) );
  LHQD1BWP \vrf/regTable_reg[7][72]  ( .E(n5105), .D(\vrf/N90 ), .Q(
        \vrf/regTable[7][72] ) );
  LHQD1BWP \vrf/regTable_reg[7][73]  ( .E(n5105), .D(\vrf/N91 ), .Q(
        \vrf/regTable[7][73] ) );
  LHQD1BWP \vrf/regTable_reg[7][74]  ( .E(n5105), .D(\vrf/N92 ), .Q(
        \vrf/regTable[7][74] ) );
  LHQD1BWP \vrf/regTable_reg[7][75]  ( .E(n5105), .D(\vrf/N93 ), .Q(
        \vrf/regTable[7][75] ) );
  LHQD1BWP \vrf/regTable_reg[7][76]  ( .E(n5105), .D(\vrf/N94 ), .Q(
        \vrf/regTable[7][76] ) );
  LHQD1BWP \vrf/regTable_reg[7][77]  ( .E(n5105), .D(\vrf/N95 ), .Q(
        \vrf/regTable[7][77] ) );
  LHQD1BWP \vrf/regTable_reg[7][78]  ( .E(n5105), .D(\vrf/N96 ), .Q(
        \vrf/regTable[7][78] ) );
  LHQD1BWP \vrf/regTable_reg[7][79]  ( .E(n5104), .D(\vrf/N97 ), .Q(
        \vrf/regTable[7][79] ) );
  LHQD1BWP \vrf/regTable_reg[7][80]  ( .E(n5104), .D(\vrf/N98 ), .Q(
        \vrf/regTable[7][80] ) );
  LHQD1BWP \vrf/regTable_reg[7][81]  ( .E(n5104), .D(\vrf/N99 ), .Q(
        \vrf/regTable[7][81] ) );
  LHQD1BWP \vrf/regTable_reg[7][82]  ( .E(n5104), .D(\vrf/N100 ), .Q(
        \vrf/regTable[7][82] ) );
  LHQD1BWP \vrf/regTable_reg[7][83]  ( .E(n5104), .D(\vrf/N101 ), .Q(
        \vrf/regTable[7][83] ) );
  LHQD1BWP \vrf/regTable_reg[7][84]  ( .E(n5104), .D(\vrf/N102 ), .Q(
        \vrf/regTable[7][84] ) );
  LHQD1BWP \vrf/regTable_reg[7][85]  ( .E(n5104), .D(\vrf/N103 ), .Q(
        \vrf/regTable[7][85] ) );
  LHQD1BWP \vrf/regTable_reg[7][86]  ( .E(n5104), .D(\vrf/N104 ), .Q(
        \vrf/regTable[7][86] ) );
  LHQD1BWP \vrf/regTable_reg[7][87]  ( .E(n5104), .D(\vrf/N105 ), .Q(
        \vrf/regTable[7][87] ) );
  LHQD1BWP \vrf/regTable_reg[7][88]  ( .E(n5104), .D(\vrf/N106 ), .Q(
        \vrf/regTable[7][88] ) );
  LHQD1BWP \vrf/regTable_reg[7][89]  ( .E(n5104), .D(\vrf/N107 ), .Q(
        \vrf/regTable[7][89] ) );
  LHQD1BWP \vrf/regTable_reg[7][90]  ( .E(n5103), .D(\vrf/N108 ), .Q(
        \vrf/regTable[7][90] ) );
  LHQD1BWP \vrf/regTable_reg[7][91]  ( .E(n5103), .D(\vrf/N109 ), .Q(
        \vrf/regTable[7][91] ) );
  LHQD1BWP \vrf/regTable_reg[7][92]  ( .E(n5103), .D(\vrf/N110 ), .Q(
        \vrf/regTable[7][92] ) );
  LHQD1BWP \vrf/regTable_reg[7][93]  ( .E(n5103), .D(\vrf/N111 ), .Q(
        \vrf/regTable[7][93] ) );
  LHQD1BWP \vrf/regTable_reg[7][94]  ( .E(n5103), .D(\vrf/N112 ), .Q(
        \vrf/regTable[7][94] ) );
  LHQD1BWP \vrf/regTable_reg[7][95]  ( .E(n5103), .D(\vrf/N113 ), .Q(
        \vrf/regTable[7][95] ) );
  LHQD1BWP \vrf/regTable_reg[7][96]  ( .E(n5103), .D(\vrf/N114 ), .Q(
        \vrf/regTable[7][96] ) );
  LHQD1BWP \vrf/regTable_reg[7][97]  ( .E(n5103), .D(\vrf/N115 ), .Q(
        \vrf/regTable[7][97] ) );
  LHQD1BWP \vrf/regTable_reg[7][98]  ( .E(n5103), .D(\vrf/N116 ), .Q(
        \vrf/regTable[7][98] ) );
  LHQD1BWP \vrf/regTable_reg[7][99]  ( .E(n5103), .D(\vrf/N118 ), .Q(
        \vrf/regTable[7][99] ) );
  LHQD1BWP \vrf/regTable_reg[7][100]  ( .E(n5113), .D(\vrf/N119 ), .Q(
        \vrf/regTable[7][100] ) );
  LHQD1BWP \vrf/regTable_reg[7][101]  ( .E(n5113), .D(\vrf/N120 ), .Q(
        \vrf/regTable[7][101] ) );
  LHQD1BWP \vrf/regTable_reg[7][102]  ( .E(n5113), .D(\vrf/N121 ), .Q(
        \vrf/regTable[7][102] ) );
  LHQD1BWP \vrf/regTable_reg[7][103]  ( .E(n5113), .D(\vrf/N122 ), .Q(
        \vrf/regTable[7][103] ) );
  LHQD1BWP \vrf/regTable_reg[7][104]  ( .E(n5113), .D(\vrf/N123 ), .Q(
        \vrf/regTable[7][104] ) );
  LHQD1BWP \vrf/regTable_reg[7][105]  ( .E(n5112), .D(\vrf/N124 ), .Q(
        \vrf/regTable[7][105] ) );
  LHQD1BWP \vrf/regTable_reg[7][106]  ( .E(n5112), .D(\vrf/N125 ), .Q(
        \vrf/regTable[7][106] ) );
  LHQD1BWP \vrf/regTable_reg[7][107]  ( .E(n5112), .D(\vrf/N126 ), .Q(
        \vrf/regTable[7][107] ) );
  LHQD1BWP \vrf/regTable_reg[7][108]  ( .E(n5112), .D(\vrf/N127 ), .Q(
        \vrf/regTable[7][108] ) );
  LHQD1BWP \vrf/regTable_reg[7][109]  ( .E(n5112), .D(\vrf/N128 ), .Q(
        \vrf/regTable[7][109] ) );
  LHQD1BWP \vrf/regTable_reg[7][110]  ( .E(n5112), .D(\vrf/N129 ), .Q(
        \vrf/regTable[7][110] ) );
  LHQD1BWP \vrf/regTable_reg[7][111]  ( .E(n5112), .D(\vrf/N130 ), .Q(
        \vrf/regTable[7][111] ) );
  LHQD1BWP \vrf/regTable_reg[7][112]  ( .E(n5112), .D(\vrf/N131 ), .Q(
        \vrf/regTable[7][112] ) );
  LHQD1BWP \vrf/regTable_reg[7][113]  ( .E(n5112), .D(\vrf/N132 ), .Q(
        \vrf/regTable[7][113] ) );
  LHQD1BWP \vrf/regTable_reg[7][114]  ( .E(n5112), .D(\vrf/N133 ), .Q(
        \vrf/regTable[7][114] ) );
  LHQD1BWP \vrf/regTable_reg[7][115]  ( .E(n5112), .D(\vrf/N134 ), .Q(
        \vrf/regTable[7][115] ) );
  LHQD1BWP \vrf/regTable_reg[7][116]  ( .E(n5111), .D(\vrf/N135 ), .Q(
        \vrf/regTable[7][116] ) );
  LHQD1BWP \vrf/regTable_reg[7][117]  ( .E(n5111), .D(\vrf/N136 ), .Q(
        \vrf/regTable[7][117] ) );
  LHQD1BWP \vrf/regTable_reg[7][118]  ( .E(n5111), .D(\vrf/N137 ), .Q(
        \vrf/regTable[7][118] ) );
  LHQD1BWP \vrf/regTable_reg[7][119]  ( .E(n5111), .D(\vrf/N138 ), .Q(
        \vrf/regTable[7][119] ) );
  LHQD1BWP \vrf/regTable_reg[7][120]  ( .E(n5111), .D(\vrf/N139 ), .Q(
        \vrf/regTable[7][120] ) );
  LHQD1BWP \vrf/regTable_reg[7][121]  ( .E(n5111), .D(\vrf/N140 ), .Q(
        \vrf/regTable[7][121] ) );
  LHQD1BWP \vrf/regTable_reg[7][122]  ( .E(n5111), .D(\vrf/N141 ), .Q(
        \vrf/regTable[7][122] ) );
  LHQD1BWP \vrf/regTable_reg[7][123]  ( .E(n5111), .D(\vrf/N142 ), .Q(
        \vrf/regTable[7][123] ) );
  LHQD1BWP \vrf/regTable_reg[7][124]  ( .E(n5111), .D(\vrf/N143 ), .Q(
        \vrf/regTable[7][124] ) );
  LHQD1BWP \vrf/regTable_reg[7][125]  ( .E(n5111), .D(\vrf/N144 ), .Q(
        \vrf/regTable[7][125] ) );
  LHQD1BWP \vrf/regTable_reg[7][126]  ( .E(n5111), .D(\vrf/N145 ), .Q(
        \vrf/regTable[7][126] ) );
  LHQD1BWP \vrf/regTable_reg[7][127]  ( .E(n5110), .D(\vrf/N146 ), .Q(
        \vrf/regTable[7][127] ) );
  LHQD1BWP \vrf/regTable_reg[7][128]  ( .E(n5113), .D(\vrf/N147 ), .Q(
        \vrf/regTable[7][128] ) );
  LHQD1BWP \vrf/regTable_reg[7][129]  ( .E(n5113), .D(\vrf/N148 ), .Q(
        \vrf/regTable[7][129] ) );
  LHQD1BWP \vrf/regTable_reg[7][130]  ( .E(n5113), .D(\vrf/N149 ), .Q(
        \vrf/regTable[7][130] ) );
  LHQD1BWP \vrf/regTable_reg[7][131]  ( .E(n5113), .D(\vrf/N150 ), .Q(
        \vrf/regTable[7][131] ) );
  LHQD1BWP \vrf/regTable_reg[7][132]  ( .E(n5113), .D(\vrf/N151 ), .Q(
        \vrf/regTable[7][132] ) );
  LHQD1BWP \vrf/regTable_reg[7][133]  ( .E(n5113), .D(\vrf/N152 ), .Q(
        \vrf/regTable[7][133] ) );
  LHQD1BWP \vrf/regTable_reg[7][134]  ( .E(n5114), .D(\vrf/N153 ), .Q(
        \vrf/regTable[7][134] ) );
  LHQD1BWP \vrf/regTable_reg[7][135]  ( .E(n5114), .D(\vrf/N154 ), .Q(
        \vrf/regTable[7][135] ) );
  LHQD1BWP \vrf/regTable_reg[7][136]  ( .E(n5114), .D(\vrf/N155 ), .Q(
        \vrf/regTable[7][136] ) );
  LHQD1BWP \vrf/regTable_reg[7][137]  ( .E(n5114), .D(\vrf/N156 ), .Q(
        \vrf/regTable[7][137] ) );
  LHQD1BWP \vrf/regTable_reg[7][138]  ( .E(n5114), .D(\vrf/N157 ), .Q(
        \vrf/regTable[7][138] ) );
  LHQD1BWP \vrf/regTable_reg[7][139]  ( .E(n5114), .D(\vrf/N158 ), .Q(
        \vrf/regTable[7][139] ) );
  LHQD1BWP \vrf/regTable_reg[7][140]  ( .E(n5114), .D(\vrf/N159 ), .Q(
        \vrf/regTable[7][140] ) );
  LHQD1BWP \vrf/regTable_reg[7][141]  ( .E(n5114), .D(\vrf/N160 ), .Q(
        \vrf/regTable[7][141] ) );
  LHQD1BWP \vrf/regTable_reg[7][142]  ( .E(n5114), .D(\vrf/N161 ), .Q(
        \vrf/regTable[7][142] ) );
  LHQD1BWP \vrf/regTable_reg[7][143]  ( .E(n5114), .D(\vrf/N162 ), .Q(
        \vrf/regTable[7][143] ) );
  LHQD1BWP \vrf/regTable_reg[7][144]  ( .E(n5114), .D(\vrf/N163 ), .Q(
        \vrf/regTable[7][144] ) );
  LHQD1BWP \vrf/regTable_reg[7][145]  ( .E(n5114), .D(\vrf/N164 ), .Q(
        \vrf/regTable[7][145] ) );
  LHQD1BWP \vrf/regTable_reg[7][146]  ( .E(n5115), .D(\vrf/N165 ), .Q(
        \vrf/regTable[7][146] ) );
  LHQD1BWP \vrf/regTable_reg[7][147]  ( .E(n5115), .D(\vrf/N166 ), .Q(
        \vrf/regTable[7][147] ) );
  LHQD1BWP \vrf/regTable_reg[7][148]  ( .E(n5115), .D(\vrf/N167 ), .Q(
        \vrf/regTable[7][148] ) );
  LHQD1BWP \vrf/regTable_reg[7][149]  ( .E(n5115), .D(\vrf/N168 ), .Q(
        \vrf/regTable[7][149] ) );
  LHQD1BWP \vrf/regTable_reg[7][150]  ( .E(n5115), .D(\vrf/N169 ), .Q(
        \vrf/regTable[7][150] ) );
  LHQD1BWP \vrf/regTable_reg[7][151]  ( .E(n5115), .D(\vrf/N170 ), .Q(
        \vrf/regTable[7][151] ) );
  LHQD1BWP \vrf/regTable_reg[7][152]  ( .E(n5115), .D(\vrf/N171 ), .Q(
        \vrf/regTable[7][152] ) );
  LHQD1BWP \vrf/regTable_reg[7][153]  ( .E(n5115), .D(\vrf/N172 ), .Q(
        \vrf/regTable[7][153] ) );
  LHQD1BWP \vrf/regTable_reg[7][154]  ( .E(n5115), .D(\vrf/N173 ), .Q(
        \vrf/regTable[7][154] ) );
  LHQD1BWP \vrf/regTable_reg[7][155]  ( .E(n5115), .D(\vrf/N174 ), .Q(
        \vrf/regTable[7][155] ) );
  LHQD1BWP \vrf/regTable_reg[7][156]  ( .E(n5115), .D(\vrf/N175 ), .Q(
        \vrf/regTable[7][156] ) );
  LHQD1BWP \vrf/regTable_reg[7][157]  ( .E(n5115), .D(\vrf/N176 ), .Q(
        \vrf/regTable[7][157] ) );
  LHQD1BWP \vrf/regTable_reg[7][158]  ( .E(n5116), .D(\vrf/N177 ), .Q(
        \vrf/regTable[7][158] ) );
  LHQD1BWP \vrf/regTable_reg[7][159]  ( .E(n5116), .D(\vrf/N178 ), .Q(
        \vrf/regTable[7][159] ) );
  LHQD1BWP \vrf/regTable_reg[7][160]  ( .E(n5116), .D(\vrf/N179 ), .Q(
        \vrf/regTable[7][160] ) );
  LHQD1BWP \vrf/regTable_reg[7][161]  ( .E(n5116), .D(\vrf/N180 ), .Q(
        \vrf/regTable[7][161] ) );
  LHQD1BWP \vrf/regTable_reg[7][162]  ( .E(n5116), .D(\vrf/N181 ), .Q(
        \vrf/regTable[7][162] ) );
  LHQD1BWP \vrf/regTable_reg[7][163]  ( .E(n5116), .D(\vrf/N182 ), .Q(
        \vrf/regTable[7][163] ) );
  LHQD1BWP \vrf/regTable_reg[7][164]  ( .E(n5116), .D(\vrf/N183 ), .Q(
        \vrf/regTable[7][164] ) );
  LHQD1BWP \vrf/regTable_reg[7][165]  ( .E(n5116), .D(\vrf/N184 ), .Q(
        \vrf/regTable[7][165] ) );
  LHQD1BWP \vrf/regTable_reg[7][166]  ( .E(n5116), .D(\vrf/N185 ), .Q(
        \vrf/regTable[7][166] ) );
  LHQD1BWP \vrf/regTable_reg[7][167]  ( .E(n5116), .D(\vrf/N186 ), .Q(
        \vrf/regTable[7][167] ) );
  LHQD1BWP \vrf/regTable_reg[7][168]  ( .E(n5116), .D(\vrf/N187 ), .Q(
        \vrf/regTable[7][168] ) );
  LHQD1BWP \vrf/regTable_reg[7][169]  ( .E(n5116), .D(\vrf/N188 ), .Q(
        \vrf/regTable[7][169] ) );
  LHQD1BWP \vrf/regTable_reg[7][170]  ( .E(n5117), .D(\vrf/N189 ), .Q(
        \vrf/regTable[7][170] ) );
  LHQD1BWP \vrf/regTable_reg[7][171]  ( .E(n5117), .D(\vrf/N190 ), .Q(
        \vrf/regTable[7][171] ) );
  LHQD1BWP \vrf/regTable_reg[7][172]  ( .E(n5117), .D(\vrf/N191 ), .Q(
        \vrf/regTable[7][172] ) );
  LHQD1BWP \vrf/regTable_reg[7][173]  ( .E(n5117), .D(\vrf/N192 ), .Q(
        \vrf/regTable[7][173] ) );
  LHQD1BWP \vrf/regTable_reg[7][174]  ( .E(n5117), .D(\vrf/N193 ), .Q(
        \vrf/regTable[7][174] ) );
  LHQD1BWP \vrf/regTable_reg[7][175]  ( .E(n5117), .D(\vrf/N194 ), .Q(
        \vrf/regTable[7][175] ) );
  LHQD1BWP \vrf/regTable_reg[7][176]  ( .E(n5117), .D(\vrf/N195 ), .Q(
        \vrf/regTable[7][176] ) );
  LHQD1BWP \vrf/regTable_reg[7][177]  ( .E(n5117), .D(\vrf/N196 ), .Q(
        \vrf/regTable[7][177] ) );
  LHQD1BWP \vrf/regTable_reg[7][178]  ( .E(n5117), .D(\vrf/N197 ), .Q(
        \vrf/regTable[7][178] ) );
  LHQD1BWP \vrf/regTable_reg[7][179]  ( .E(n5117), .D(\vrf/N198 ), .Q(
        \vrf/regTable[7][179] ) );
  LHQD1BWP \vrf/regTable_reg[7][180]  ( .E(n5117), .D(\vrf/N199 ), .Q(
        \vrf/regTable[7][180] ) );
  LHQD1BWP \vrf/regTable_reg[7][181]  ( .E(n5117), .D(\vrf/N200 ), .Q(
        \vrf/regTable[7][181] ) );
  LHQD1BWP \vrf/regTable_reg[7][182]  ( .E(n5118), .D(\vrf/N201 ), .Q(
        \vrf/regTable[7][182] ) );
  LHQD1BWP \vrf/regTable_reg[7][183]  ( .E(n5118), .D(\vrf/N202 ), .Q(
        \vrf/regTable[7][183] ) );
  LHQD1BWP \vrf/regTable_reg[7][184]  ( .E(n5118), .D(\vrf/N203 ), .Q(
        \vrf/regTable[7][184] ) );
  LHQD1BWP \vrf/regTable_reg[7][185]  ( .E(n5118), .D(\vrf/N204 ), .Q(
        \vrf/regTable[7][185] ) );
  LHQD1BWP \vrf/regTable_reg[7][186]  ( .E(n5118), .D(\vrf/N205 ), .Q(
        \vrf/regTable[7][186] ) );
  LHQD1BWP \vrf/regTable_reg[7][187]  ( .E(n5118), .D(\vrf/N206 ), .Q(
        \vrf/regTable[7][187] ) );
  LHQD1BWP \vrf/regTable_reg[7][188]  ( .E(n5118), .D(\vrf/N207 ), .Q(
        \vrf/regTable[7][188] ) );
  LHQD1BWP \vrf/regTable_reg[7][189]  ( .E(n5118), .D(\vrf/N208 ), .Q(
        \vrf/regTable[7][189] ) );
  LHQD1BWP \vrf/regTable_reg[7][190]  ( .E(n5118), .D(\vrf/N209 ), .Q(
        \vrf/regTable[7][190] ) );
  LHQD1BWP \vrf/regTable_reg[7][191]  ( .E(n5118), .D(\vrf/N210 ), .Q(
        \vrf/regTable[7][191] ) );
  LHQD1BWP \vrf/regTable_reg[7][192]  ( .E(n5118), .D(\vrf/N211 ), .Q(
        \vrf/regTable[7][192] ) );
  LHQD1BWP \vrf/regTable_reg[7][193]  ( .E(n5118), .D(\vrf/N212 ), .Q(
        \vrf/regTable[7][193] ) );
  LHQD1BWP \vrf/regTable_reg[7][194]  ( .E(n5119), .D(\vrf/N213 ), .Q(
        \vrf/regTable[7][194] ) );
  LHQD1BWP \vrf/regTable_reg[7][195]  ( .E(n5119), .D(\vrf/N214 ), .Q(
        \vrf/regTable[7][195] ) );
  LHQD1BWP \vrf/regTable_reg[7][196]  ( .E(n5119), .D(\vrf/N215 ), .Q(
        \vrf/regTable[7][196] ) );
  LHQD1BWP \vrf/regTable_reg[7][197]  ( .E(n5119), .D(\vrf/N216 ), .Q(
        \vrf/regTable[7][197] ) );
  LHQD1BWP \vrf/regTable_reg[7][198]  ( .E(n5119), .D(\vrf/N218 ), .Q(
        \vrf/regTable[7][198] ) );
  LHQD1BWP \vrf/regTable_reg[7][199]  ( .E(n5119), .D(\vrf/N219 ), .Q(
        \vrf/regTable[7][199] ) );
  LHQD1BWP \vrf/regTable_reg[7][200]  ( .E(n5119), .D(\vrf/N220 ), .Q(
        \vrf/regTable[7][200] ) );
  LHQD1BWP \vrf/regTable_reg[7][201]  ( .E(n5119), .D(\vrf/N221 ), .Q(
        \vrf/regTable[7][201] ) );
  LHQD1BWP \vrf/regTable_reg[7][202]  ( .E(n5119), .D(\vrf/N222 ), .Q(
        \vrf/regTable[7][202] ) );
  LHQD1BWP \vrf/regTable_reg[7][203]  ( .E(n5119), .D(\vrf/N223 ), .Q(
        \vrf/regTable[7][203] ) );
  LHQD1BWP \vrf/regTable_reg[7][204]  ( .E(n5119), .D(\vrf/N224 ), .Q(
        \vrf/regTable[7][204] ) );
  LHQD1BWP \vrf/regTable_reg[7][205]  ( .E(n5119), .D(\vrf/N225 ), .Q(
        \vrf/regTable[7][205] ) );
  LHQD1BWP \vrf/regTable_reg[7][206]  ( .E(n5120), .D(\vrf/N226 ), .Q(
        \vrf/regTable[7][206] ) );
  LHQD1BWP \vrf/regTable_reg[7][207]  ( .E(n5120), .D(\vrf/N227 ), .Q(
        \vrf/regTable[7][207] ) );
  LHQD1BWP \vrf/regTable_reg[7][208]  ( .E(n5120), .D(\vrf/N228 ), .Q(
        \vrf/regTable[7][208] ) );
  LHQD1BWP \vrf/regTable_reg[7][209]  ( .E(n5120), .D(\vrf/N229 ), .Q(
        \vrf/regTable[7][209] ) );
  LHQD1BWP \vrf/regTable_reg[7][210]  ( .E(n5120), .D(\vrf/N230 ), .Q(
        \vrf/regTable[7][210] ) );
  LHQD1BWP \vrf/regTable_reg[7][211]  ( .E(n5120), .D(\vrf/N231 ), .Q(
        \vrf/regTable[7][211] ) );
  LHQD1BWP \vrf/regTable_reg[7][212]  ( .E(n5120), .D(\vrf/N232 ), .Q(
        \vrf/regTable[7][212] ) );
  LHQD1BWP \vrf/regTable_reg[7][213]  ( .E(n5120), .D(\vrf/N233 ), .Q(
        \vrf/regTable[7][213] ) );
  LHQD1BWP \vrf/regTable_reg[7][214]  ( .E(n5120), .D(\vrf/N234 ), .Q(
        \vrf/regTable[7][214] ) );
  LHQD1BWP \vrf/regTable_reg[7][215]  ( .E(n5120), .D(\vrf/N235 ), .Q(
        \vrf/regTable[7][215] ) );
  LHQD1BWP \vrf/regTable_reg[7][216]  ( .E(n5120), .D(\vrf/N236 ), .Q(
        \vrf/regTable[7][216] ) );
  LHQD1BWP \vrf/regTable_reg[7][217]  ( .E(n5120), .D(\vrf/N237 ), .Q(
        \vrf/regTable[7][217] ) );
  LHQD1BWP \vrf/regTable_reg[7][218]  ( .E(n5121), .D(\vrf/N238 ), .Q(
        \vrf/regTable[7][218] ) );
  LHQD1BWP \vrf/regTable_reg[7][219]  ( .E(n5121), .D(\vrf/N239 ), .Q(
        \vrf/regTable[7][219] ) );
  LHQD1BWP \vrf/regTable_reg[7][220]  ( .E(n5121), .D(\vrf/N240 ), .Q(
        \vrf/regTable[7][220] ) );
  LHQD1BWP \vrf/regTable_reg[7][221]  ( .E(n5121), .D(\vrf/N241 ), .Q(
        \vrf/regTable[7][221] ) );
  LHQD1BWP \vrf/regTable_reg[7][222]  ( .E(n5121), .D(\vrf/N242 ), .Q(
        \vrf/regTable[7][222] ) );
  LHQD1BWP \vrf/regTable_reg[7][223]  ( .E(n5121), .D(\vrf/N243 ), .Q(
        \vrf/regTable[7][223] ) );
  LHQD1BWP \vrf/regTable_reg[7][224]  ( .E(n5121), .D(\vrf/N244 ), .Q(
        \vrf/regTable[7][224] ) );
  LHQD1BWP \vrf/regTable_reg[7][225]  ( .E(n5121), .D(\vrf/N245 ), .Q(
        \vrf/regTable[7][225] ) );
  LHQD1BWP \vrf/regTable_reg[7][226]  ( .E(n5121), .D(\vrf/N246 ), .Q(
        \vrf/regTable[7][226] ) );
  LHQD1BWP \vrf/regTable_reg[7][227]  ( .E(n5121), .D(\vrf/N247 ), .Q(
        \vrf/regTable[7][227] ) );
  LHQD1BWP \vrf/regTable_reg[7][228]  ( .E(n5121), .D(\vrf/N248 ), .Q(
        \vrf/regTable[7][228] ) );
  LHQD1BWP \vrf/regTable_reg[7][229]  ( .E(n5121), .D(\vrf/N249 ), .Q(
        \vrf/regTable[7][229] ) );
  LHQD1BWP \vrf/regTable_reg[7][230]  ( .E(n5122), .D(\vrf/N250 ), .Q(
        \vrf/regTable[7][230] ) );
  LHQD1BWP \vrf/regTable_reg[7][231]  ( .E(n5122), .D(\vrf/N251 ), .Q(
        \vrf/regTable[7][231] ) );
  LHQD1BWP \vrf/regTable_reg[7][232]  ( .E(n5122), .D(\vrf/N252 ), .Q(
        \vrf/regTable[7][232] ) );
  LHQD1BWP \vrf/regTable_reg[7][233]  ( .E(n5122), .D(\vrf/N253 ), .Q(
        \vrf/regTable[7][233] ) );
  LHQD1BWP \vrf/regTable_reg[7][234]  ( .E(n5122), .D(\vrf/N254 ), .Q(
        \vrf/regTable[7][234] ) );
  LHQD1BWP \vrf/regTable_reg[7][235]  ( .E(n5122), .D(\vrf/N255 ), .Q(
        \vrf/regTable[7][235] ) );
  LHQD1BWP \vrf/regTable_reg[7][236]  ( .E(n5122), .D(\vrf/N256 ), .Q(
        \vrf/regTable[7][236] ) );
  LHQD1BWP \vrf/regTable_reg[7][237]  ( .E(n5122), .D(\vrf/N257 ), .Q(
        \vrf/regTable[7][237] ) );
  LHQD1BWP \vrf/regTable_reg[7][238]  ( .E(n5122), .D(\vrf/N258 ), .Q(
        \vrf/regTable[7][238] ) );
  LHQD1BWP \vrf/regTable_reg[7][239]  ( .E(n5122), .D(\vrf/N259 ), .Q(
        \vrf/regTable[7][239] ) );
  LHQD1BWP \vrf/regTable_reg[7][240]  ( .E(n5122), .D(\vrf/N260 ), .Q(
        \vrf/regTable[7][240] ) );
  LHQD1BWP \vrf/regTable_reg[7][241]  ( .E(n5122), .D(\vrf/N261 ), .Q(
        \vrf/regTable[7][241] ) );
  LHQD1BWP \vrf/regTable_reg[7][242]  ( .E(n5123), .D(\vrf/N262 ), .Q(
        \vrf/regTable[7][242] ) );
  LHQD1BWP \vrf/regTable_reg[7][243]  ( .E(n5123), .D(\vrf/N263 ), .Q(
        \vrf/regTable[7][243] ) );
  LHQD1BWP \vrf/regTable_reg[7][244]  ( .E(n5123), .D(\vrf/N264 ), .Q(
        \vrf/regTable[7][244] ) );
  LHQD1BWP \vrf/regTable_reg[7][245]  ( .E(n5123), .D(\vrf/N265 ), .Q(
        \vrf/regTable[7][245] ) );
  LHQD1BWP \vrf/regTable_reg[7][246]  ( .E(n5123), .D(\vrf/N266 ), .Q(
        \vrf/regTable[7][246] ) );
  LHQD1BWP \vrf/regTable_reg[7][247]  ( .E(n5123), .D(\vrf/N267 ), .Q(
        \vrf/regTable[7][247] ) );
  LHQD1BWP \vrf/regTable_reg[7][248]  ( .E(n5123), .D(\vrf/N268 ), .Q(
        \vrf/regTable[7][248] ) );
  LHQD1BWP \vrf/regTable_reg[7][249]  ( .E(n5123), .D(\vrf/N269 ), .Q(
        \vrf/regTable[7][249] ) );
  LHQD1BWP \vrf/regTable_reg[7][250]  ( .E(n5123), .D(\vrf/N270 ), .Q(
        \vrf/regTable[7][250] ) );
  LHQD1BWP \vrf/regTable_reg[7][251]  ( .E(n5123), .D(\vrf/N271 ), .Q(
        \vrf/regTable[7][251] ) );
  LHQD1BWP \vrf/regTable_reg[7][252]  ( .E(n5123), .D(\vrf/N272 ), .Q(
        \vrf/regTable[7][252] ) );
  LHQD1BWP \vrf/regTable_reg[7][253]  ( .E(n5123), .D(\vrf/N273 ), .Q(
        \vrf/regTable[7][253] ) );
  LHQD1BWP \vrf/regTable_reg[3][0]  ( .E(n5249), .D(\vrf/N18 ), .Q(
        \vrf/regTable[3][0] ) );
  LHQD1BWP \vrf/regTable_reg[3][1]  ( .E(n5246), .D(\vrf/N19 ), .Q(
        \vrf/regTable[3][1] ) );
  LHQD1BWP \vrf/regTable_reg[3][2]  ( .E(n5245), .D(\vrf/N20 ), .Q(
        \vrf/regTable[3][2] ) );
  LHQD1BWP \vrf/regTable_reg[3][3]  ( .E(n5244), .D(\vrf/N21 ), .Q(
        \vrf/regTable[3][3] ) );
  LHQD1BWP \vrf/regTable_reg[3][4]  ( .E(n5243), .D(\vrf/N22 ), .Q(
        \vrf/regTable[3][4] ) );
  LHQD1BWP \vrf/regTable_reg[3][5]  ( .E(n5242), .D(\vrf/N23 ), .Q(
        \vrf/regTable[3][5] ) );
  LHQD1BWP \vrf/regTable_reg[3][6]  ( .E(n5241), .D(\vrf/N24 ), .Q(
        \vrf/regTable[3][6] ) );
  LHQD1BWP \vrf/regTable_reg[3][7]  ( .E(n5240), .D(\vrf/N25 ), .Q(
        \vrf/regTable[3][7] ) );
  LHQD1BWP \vrf/regTable_reg[3][8]  ( .E(n5239), .D(\vrf/N26 ), .Q(
        \vrf/regTable[3][8] ) );
  LHQD1BWP \vrf/regTable_reg[3][9]  ( .E(n5239), .D(\vrf/N27 ), .Q(
        \vrf/regTable[3][9] ) );
  LHQD1BWP \vrf/regTable_reg[3][10]  ( .E(n5248), .D(\vrf/N28 ), .Q(
        \vrf/regTable[3][10] ) );
  LHQD1BWP \vrf/regTable_reg[3][11]  ( .E(n5247), .D(\vrf/N29 ), .Q(
        \vrf/regTable[3][11] ) );
  LHQD1BWP \vrf/regTable_reg[3][12]  ( .E(n5246), .D(\vrf/N30 ), .Q(
        \vrf/regTable[3][12] ) );
  LHQD1BWP \vrf/regTable_reg[3][13]  ( .E(n5246), .D(\vrf/N31 ), .Q(
        \vrf/regTable[3][13] ) );
  LHQD1BWP \vrf/regTable_reg[3][14]  ( .E(n5246), .D(\vrf/N32 ), .Q(
        \vrf/regTable[3][14] ) );
  LHQD1BWP \vrf/regTable_reg[3][17]  ( .E(n5246), .D(\vrf/N35 ), .Q(
        \vrf/regTable[3][17] ) );
  LHQD1BWP \vrf/regTable_reg[3][18]  ( .E(n5246), .D(\vrf/N36 ), .Q(
        \vrf/regTable[3][18] ) );
  LHQD1BWP \vrf/regTable_reg[3][19]  ( .E(n5246), .D(\vrf/N37 ), .Q(
        \vrf/regTable[3][19] ) );
  LHQD1BWP \vrf/regTable_reg[3][20]  ( .E(n5246), .D(\vrf/N38 ), .Q(
        \vrf/regTable[3][20] ) );
  LHQD1BWP \vrf/regTable_reg[3][21]  ( .E(n5246), .D(\vrf/N39 ), .Q(
        \vrf/regTable[3][21] ) );
  LHQD1BWP \vrf/regTable_reg[3][22]  ( .E(n5246), .D(\vrf/N40 ), .Q(
        \vrf/regTable[3][22] ) );
  LHQD1BWP \vrf/regTable_reg[3][23]  ( .E(n5246), .D(\vrf/N41 ), .Q(
        \vrf/regTable[3][23] ) );
  LHQD1BWP \vrf/regTable_reg[3][24]  ( .E(n5245), .D(\vrf/N42 ), .Q(
        \vrf/regTable[3][24] ) );
  LHQD1BWP \vrf/regTable_reg[3][25]  ( .E(n5245), .D(\vrf/N43 ), .Q(
        \vrf/regTable[3][25] ) );
  LHQD1BWP \vrf/regTable_reg[3][26]  ( .E(n5245), .D(\vrf/N44 ), .Q(
        \vrf/regTable[3][26] ) );
  LHQD1BWP \vrf/regTable_reg[3][27]  ( .E(n5245), .D(\vrf/N45 ), .Q(
        \vrf/regTable[3][27] ) );
  LHQD1BWP \vrf/regTable_reg[3][28]  ( .E(n5245), .D(\vrf/N46 ), .Q(
        \vrf/regTable[3][28] ) );
  LHQD1BWP \vrf/regTable_reg[3][29]  ( .E(n5245), .D(\vrf/N47 ), .Q(
        \vrf/regTable[3][29] ) );
  LHQD1BWP \vrf/regTable_reg[3][30]  ( .E(n5245), .D(\vrf/N48 ), .Q(
        \vrf/regTable[3][30] ) );
  LHQD1BWP \vrf/regTable_reg[3][31]  ( .E(n5245), .D(\vrf/N49 ), .Q(
        \vrf/regTable[3][31] ) );
  LHQD1BWP \vrf/regTable_reg[3][32]  ( .E(n5245), .D(\vrf/N50 ), .Q(
        \vrf/regTable[3][32] ) );
  LHQD1BWP \vrf/regTable_reg[3][33]  ( .E(n5245), .D(\vrf/N51 ), .Q(
        \vrf/regTable[3][33] ) );
  LHQD1BWP \vrf/regTable_reg[3][34]  ( .E(n5245), .D(\vrf/N52 ), .Q(
        \vrf/regTable[3][34] ) );
  LHQD1BWP \vrf/regTable_reg[3][35]  ( .E(n5244), .D(\vrf/N53 ), .Q(
        \vrf/regTable[3][35] ) );
  LHQD1BWP \vrf/regTable_reg[3][36]  ( .E(n5244), .D(\vrf/N54 ), .Q(
        \vrf/regTable[3][36] ) );
  LHQD1BWP \vrf/regTable_reg[3][37]  ( .E(n5244), .D(\vrf/N55 ), .Q(
        \vrf/regTable[3][37] ) );
  LHQD1BWP \vrf/regTable_reg[3][38]  ( .E(n5244), .D(\vrf/N56 ), .Q(
        \vrf/regTable[3][38] ) );
  LHQD1BWP \vrf/regTable_reg[3][39]  ( .E(n5244), .D(\vrf/N57 ), .Q(
        \vrf/regTable[3][39] ) );
  LHQD1BWP \vrf/regTable_reg[3][40]  ( .E(n5244), .D(\vrf/N58 ), .Q(
        \vrf/regTable[3][40] ) );
  LHQD1BWP \vrf/regTable_reg[3][41]  ( .E(n5244), .D(\vrf/N59 ), .Q(
        \vrf/regTable[3][41] ) );
  LHQD1BWP \vrf/regTable_reg[3][42]  ( .E(n5244), .D(\vrf/N60 ), .Q(
        \vrf/regTable[3][42] ) );
  LHQD1BWP \vrf/regTable_reg[3][43]  ( .E(n5244), .D(\vrf/N61 ), .Q(
        \vrf/regTable[3][43] ) );
  LHQD1BWP \vrf/regTable_reg[3][44]  ( .E(n5244), .D(\vrf/N62 ), .Q(
        \vrf/regTable[3][44] ) );
  LHQD1BWP \vrf/regTable_reg[3][45]  ( .E(n5244), .D(\vrf/N63 ), .Q(
        \vrf/regTable[3][45] ) );
  LHQD1BWP \vrf/regTable_reg[3][46]  ( .E(n5243), .D(\vrf/N64 ), .Q(
        \vrf/regTable[3][46] ) );
  LHQD1BWP \vrf/regTable_reg[3][47]  ( .E(n5243), .D(\vrf/N65 ), .Q(
        \vrf/regTable[3][47] ) );
  LHQD1BWP \vrf/regTable_reg[3][48]  ( .E(n5243), .D(\vrf/N66 ), .Q(
        \vrf/regTable[3][48] ) );
  LHQD1BWP \vrf/regTable_reg[3][49]  ( .E(n5243), .D(\vrf/N67 ), .Q(
        \vrf/regTable[3][49] ) );
  LHQD1BWP \vrf/regTable_reg[3][50]  ( .E(n5243), .D(\vrf/N68 ), .Q(
        \vrf/regTable[3][50] ) );
  LHQD1BWP \vrf/regTable_reg[3][51]  ( .E(n5243), .D(\vrf/N69 ), .Q(
        \vrf/regTable[3][51] ) );
  LHQD1BWP \vrf/regTable_reg[3][52]  ( .E(n5243), .D(\vrf/N70 ), .Q(
        \vrf/regTable[3][52] ) );
  LHQD1BWP \vrf/regTable_reg[3][53]  ( .E(n5243), .D(\vrf/N71 ), .Q(
        \vrf/regTable[3][53] ) );
  LHQD1BWP \vrf/regTable_reg[3][54]  ( .E(n5243), .D(\vrf/N72 ), .Q(
        \vrf/regTable[3][54] ) );
  LHQD1BWP \vrf/regTable_reg[3][55]  ( .E(n5243), .D(\vrf/N73 ), .Q(
        \vrf/regTable[3][55] ) );
  LHQD1BWP \vrf/regTable_reg[3][56]  ( .E(n5243), .D(\vrf/N74 ), .Q(
        \vrf/regTable[3][56] ) );
  LHQD1BWP \vrf/regTable_reg[3][57]  ( .E(n5242), .D(\vrf/N75 ), .Q(
        \vrf/regTable[3][57] ) );
  LHQD1BWP \vrf/regTable_reg[3][58]  ( .E(n5242), .D(\vrf/N76 ), .Q(
        \vrf/regTable[3][58] ) );
  LHQD1BWP \vrf/regTable_reg[3][59]  ( .E(n5242), .D(\vrf/N77 ), .Q(
        \vrf/regTable[3][59] ) );
  LHQD1BWP \vrf/regTable_reg[3][60]  ( .E(n5242), .D(\vrf/N78 ), .Q(
        \vrf/regTable[3][60] ) );
  LHQD1BWP \vrf/regTable_reg[3][61]  ( .E(n5242), .D(\vrf/N79 ), .Q(
        \vrf/regTable[3][61] ) );
  LHQD1BWP \vrf/regTable_reg[3][62]  ( .E(n5242), .D(\vrf/N80 ), .Q(
        \vrf/regTable[3][62] ) );
  LHQD1BWP \vrf/regTable_reg[3][63]  ( .E(n5242), .D(\vrf/N81 ), .Q(
        \vrf/regTable[3][63] ) );
  LHQD1BWP \vrf/regTable_reg[3][64]  ( .E(n5242), .D(\vrf/N82 ), .Q(
        \vrf/regTable[3][64] ) );
  LHQD1BWP \vrf/regTable_reg[3][65]  ( .E(n5242), .D(\vrf/N83 ), .Q(
        \vrf/regTable[3][65] ) );
  LHQD1BWP \vrf/regTable_reg[3][66]  ( .E(n5242), .D(\vrf/N84 ), .Q(
        \vrf/regTable[3][66] ) );
  LHQD1BWP \vrf/regTable_reg[3][67]  ( .E(n5242), .D(\vrf/N85 ), .Q(
        \vrf/regTable[3][67] ) );
  LHQD1BWP \vrf/regTable_reg[3][68]  ( .E(n5241), .D(\vrf/N86 ), .Q(
        \vrf/regTable[3][68] ) );
  LHQD1BWP \vrf/regTable_reg[3][69]  ( .E(n5241), .D(\vrf/N87 ), .Q(
        \vrf/regTable[3][69] ) );
  LHQD1BWP \vrf/regTable_reg[3][70]  ( .E(n5241), .D(\vrf/N88 ), .Q(
        \vrf/regTable[3][70] ) );
  LHQD1BWP \vrf/regTable_reg[3][71]  ( .E(n5241), .D(\vrf/N89 ), .Q(
        \vrf/regTable[3][71] ) );
  LHQD1BWP \vrf/regTable_reg[3][72]  ( .E(n5241), .D(\vrf/N90 ), .Q(
        \vrf/regTable[3][72] ) );
  LHQD1BWP \vrf/regTable_reg[3][73]  ( .E(n5241), .D(\vrf/N91 ), .Q(
        \vrf/regTable[3][73] ) );
  LHQD1BWP \vrf/regTable_reg[3][74]  ( .E(n5241), .D(\vrf/N92 ), .Q(
        \vrf/regTable[3][74] ) );
  LHQD1BWP \vrf/regTable_reg[3][75]  ( .E(n5241), .D(\vrf/N93 ), .Q(
        \vrf/regTable[3][75] ) );
  LHQD1BWP \vrf/regTable_reg[3][76]  ( .E(n5241), .D(\vrf/N94 ), .Q(
        \vrf/regTable[3][76] ) );
  LHQD1BWP \vrf/regTable_reg[3][77]  ( .E(n5241), .D(\vrf/N95 ), .Q(
        \vrf/regTable[3][77] ) );
  LHQD1BWP \vrf/regTable_reg[3][78]  ( .E(n5241), .D(\vrf/N96 ), .Q(
        \vrf/regTable[3][78] ) );
  LHQD1BWP \vrf/regTable_reg[3][79]  ( .E(n5240), .D(\vrf/N97 ), .Q(
        \vrf/regTable[3][79] ) );
  LHQD1BWP \vrf/regTable_reg[3][80]  ( .E(n5240), .D(\vrf/N98 ), .Q(
        \vrf/regTable[3][80] ) );
  LHQD1BWP \vrf/regTable_reg[3][81]  ( .E(n5240), .D(\vrf/N99 ), .Q(
        \vrf/regTable[3][81] ) );
  LHQD1BWP \vrf/regTable_reg[3][82]  ( .E(n5240), .D(\vrf/N100 ), .Q(
        \vrf/regTable[3][82] ) );
  LHQD1BWP \vrf/regTable_reg[3][83]  ( .E(n5240), .D(\vrf/N101 ), .Q(
        \vrf/regTable[3][83] ) );
  LHQD1BWP \vrf/regTable_reg[3][84]  ( .E(n5240), .D(\vrf/N102 ), .Q(
        \vrf/regTable[3][84] ) );
  LHQD1BWP \vrf/regTable_reg[3][85]  ( .E(n5240), .D(\vrf/N103 ), .Q(
        \vrf/regTable[3][85] ) );
  LHQD1BWP \vrf/regTable_reg[3][86]  ( .E(n5240), .D(\vrf/N104 ), .Q(
        \vrf/regTable[3][86] ) );
  LHQD1BWP \vrf/regTable_reg[3][87]  ( .E(n5240), .D(\vrf/N105 ), .Q(
        \vrf/regTable[3][87] ) );
  LHQD1BWP \vrf/regTable_reg[3][88]  ( .E(n5240), .D(\vrf/N106 ), .Q(
        \vrf/regTable[3][88] ) );
  LHQD1BWP \vrf/regTable_reg[3][89]  ( .E(n5240), .D(\vrf/N107 ), .Q(
        \vrf/regTable[3][89] ) );
  LHQD1BWP \vrf/regTable_reg[3][90]  ( .E(n5239), .D(\vrf/N108 ), .Q(
        \vrf/regTable[3][90] ) );
  LHQD1BWP \vrf/regTable_reg[3][91]  ( .E(n5239), .D(\vrf/N109 ), .Q(
        \vrf/regTable[3][91] ) );
  LHQD1BWP \vrf/regTable_reg[3][92]  ( .E(n5239), .D(\vrf/N110 ), .Q(
        \vrf/regTable[3][92] ) );
  LHQD1BWP \vrf/regTable_reg[3][93]  ( .E(n5239), .D(\vrf/N111 ), .Q(
        \vrf/regTable[3][93] ) );
  LHQD1BWP \vrf/regTable_reg[3][94]  ( .E(n5239), .D(\vrf/N112 ), .Q(
        \vrf/regTable[3][94] ) );
  LHQD1BWP \vrf/regTable_reg[3][95]  ( .E(n5239), .D(\vrf/N113 ), .Q(
        \vrf/regTable[3][95] ) );
  LHQD1BWP \vrf/regTable_reg[3][96]  ( .E(n5239), .D(\vrf/N114 ), .Q(
        \vrf/regTable[3][96] ) );
  LHQD1BWP \vrf/regTable_reg[3][97]  ( .E(n5239), .D(\vrf/N115 ), .Q(
        \vrf/regTable[3][97] ) );
  LHQD1BWP \vrf/regTable_reg[3][98]  ( .E(n5239), .D(\vrf/N116 ), .Q(
        \vrf/regTable[3][98] ) );
  LHQD1BWP \vrf/regTable_reg[3][99]  ( .E(n5239), .D(\vrf/N118 ), .Q(
        \vrf/regTable[3][99] ) );
  LHQD1BWP \vrf/regTable_reg[3][100]  ( .E(n5249), .D(\vrf/N119 ), .Q(
        \vrf/regTable[3][100] ) );
  LHQD1BWP \vrf/regTable_reg[3][101]  ( .E(n5249), .D(\vrf/N120 ), .Q(
        \vrf/regTable[3][101] ) );
  LHQD1BWP \vrf/regTable_reg[3][102]  ( .E(n5249), .D(\vrf/N121 ), .Q(
        \vrf/regTable[3][102] ) );
  LHQD1BWP \vrf/regTable_reg[3][103]  ( .E(n5249), .D(\vrf/N122 ), .Q(
        \vrf/regTable[3][103] ) );
  LHQD1BWP \vrf/regTable_reg[3][104]  ( .E(n5249), .D(\vrf/N123 ), .Q(
        \vrf/regTable[3][104] ) );
  LHQD1BWP \vrf/regTable_reg[3][105]  ( .E(n5248), .D(\vrf/N124 ), .Q(
        \vrf/regTable[3][105] ) );
  LHQD1BWP \vrf/regTable_reg[3][106]  ( .E(n5248), .D(\vrf/N125 ), .Q(
        \vrf/regTable[3][106] ) );
  LHQD1BWP \vrf/regTable_reg[3][107]  ( .E(n5248), .D(\vrf/N126 ), .Q(
        \vrf/regTable[3][107] ) );
  LHQD1BWP \vrf/regTable_reg[3][108]  ( .E(n5248), .D(\vrf/N127 ), .Q(
        \vrf/regTable[3][108] ) );
  LHQD1BWP \vrf/regTable_reg[3][109]  ( .E(n5248), .D(\vrf/N128 ), .Q(
        \vrf/regTable[3][109] ) );
  LHQD1BWP \vrf/regTable_reg[3][110]  ( .E(n5248), .D(\vrf/N129 ), .Q(
        \vrf/regTable[3][110] ) );
  LHQD1BWP \vrf/regTable_reg[3][111]  ( .E(n5248), .D(\vrf/N130 ), .Q(
        \vrf/regTable[3][111] ) );
  LHQD1BWP \vrf/regTable_reg[3][112]  ( .E(n5248), .D(\vrf/N131 ), .Q(
        \vrf/regTable[3][112] ) );
  LHQD1BWP \vrf/regTable_reg[3][113]  ( .E(n5248), .D(\vrf/N132 ), .Q(
        \vrf/regTable[3][113] ) );
  LHQD1BWP \vrf/regTable_reg[3][114]  ( .E(n5248), .D(\vrf/N133 ), .Q(
        \vrf/regTable[3][114] ) );
  LHQD1BWP \vrf/regTable_reg[3][115]  ( .E(n5248), .D(\vrf/N134 ), .Q(
        \vrf/regTable[3][115] ) );
  LHQD1BWP \vrf/regTable_reg[3][116]  ( .E(n5247), .D(\vrf/N135 ), .Q(
        \vrf/regTable[3][116] ) );
  LHQD1BWP \vrf/regTable_reg[3][117]  ( .E(n5247), .D(\vrf/N136 ), .Q(
        \vrf/regTable[3][117] ) );
  LHQD1BWP \vrf/regTable_reg[3][118]  ( .E(n5247), .D(\vrf/N137 ), .Q(
        \vrf/regTable[3][118] ) );
  LHQD1BWP \vrf/regTable_reg[3][119]  ( .E(n5247), .D(\vrf/N138 ), .Q(
        \vrf/regTable[3][119] ) );
  LHQD1BWP \vrf/regTable_reg[3][120]  ( .E(n5247), .D(\vrf/N139 ), .Q(
        \vrf/regTable[3][120] ) );
  LHQD1BWP \vrf/regTable_reg[3][121]  ( .E(n5247), .D(\vrf/N140 ), .Q(
        \vrf/regTable[3][121] ) );
  LHQD1BWP \vrf/regTable_reg[3][122]  ( .E(n5247), .D(\vrf/N141 ), .Q(
        \vrf/regTable[3][122] ) );
  LHQD1BWP \vrf/regTable_reg[3][123]  ( .E(n5247), .D(\vrf/N142 ), .Q(
        \vrf/regTable[3][123] ) );
  LHQD1BWP \vrf/regTable_reg[3][124]  ( .E(n5247), .D(\vrf/N143 ), .Q(
        \vrf/regTable[3][124] ) );
  LHQD1BWP \vrf/regTable_reg[3][125]  ( .E(n5247), .D(\vrf/N144 ), .Q(
        \vrf/regTable[3][125] ) );
  LHQD1BWP \vrf/regTable_reg[3][126]  ( .E(n5247), .D(\vrf/N145 ), .Q(
        \vrf/regTable[3][126] ) );
  LHQD1BWP \vrf/regTable_reg[3][127]  ( .E(n5246), .D(\vrf/N146 ), .Q(
        \vrf/regTable[3][127] ) );
  LHQD1BWP \vrf/regTable_reg[3][128]  ( .E(n5249), .D(\vrf/N147 ), .Q(
        \vrf/regTable[3][128] ) );
  LHQD1BWP \vrf/regTable_reg[3][129]  ( .E(n5249), .D(\vrf/N148 ), .Q(
        \vrf/regTable[3][129] ) );
  LHQD1BWP \vrf/regTable_reg[3][130]  ( .E(n5249), .D(\vrf/N149 ), .Q(
        \vrf/regTable[3][130] ) );
  LHQD1BWP \vrf/regTable_reg[3][131]  ( .E(n5249), .D(\vrf/N150 ), .Q(
        \vrf/regTable[3][131] ) );
  LHQD1BWP \vrf/regTable_reg[3][132]  ( .E(n5249), .D(\vrf/N151 ), .Q(
        \vrf/regTable[3][132] ) );
  LHQD1BWP \vrf/regTable_reg[3][133]  ( .E(n5249), .D(\vrf/N152 ), .Q(
        \vrf/regTable[3][133] ) );
  LHQD1BWP \vrf/regTable_reg[3][134]  ( .E(n5250), .D(\vrf/N153 ), .Q(
        \vrf/regTable[3][134] ) );
  LHQD1BWP \vrf/regTable_reg[3][135]  ( .E(n5250), .D(\vrf/N154 ), .Q(
        \vrf/regTable[3][135] ) );
  LHQD1BWP \vrf/regTable_reg[3][136]  ( .E(n5250), .D(\vrf/N155 ), .Q(
        \vrf/regTable[3][136] ) );
  LHQD1BWP \vrf/regTable_reg[3][137]  ( .E(n5250), .D(\vrf/N156 ), .Q(
        \vrf/regTable[3][137] ) );
  LHQD1BWP \vrf/regTable_reg[3][138]  ( .E(n5250), .D(\vrf/N157 ), .Q(
        \vrf/regTable[3][138] ) );
  LHQD1BWP \vrf/regTable_reg[3][139]  ( .E(n5250), .D(\vrf/N158 ), .Q(
        \vrf/regTable[3][139] ) );
  LHQD1BWP \vrf/regTable_reg[3][140]  ( .E(n5250), .D(\vrf/N159 ), .Q(
        \vrf/regTable[3][140] ) );
  LHQD1BWP \vrf/regTable_reg[3][141]  ( .E(n5250), .D(\vrf/N160 ), .Q(
        \vrf/regTable[3][141] ) );
  LHQD1BWP \vrf/regTable_reg[3][142]  ( .E(n5250), .D(\vrf/N161 ), .Q(
        \vrf/regTable[3][142] ) );
  LHQD1BWP \vrf/regTable_reg[3][143]  ( .E(n5250), .D(\vrf/N162 ), .Q(
        \vrf/regTable[3][143] ) );
  LHQD1BWP \vrf/regTable_reg[3][144]  ( .E(n5250), .D(\vrf/N163 ), .Q(
        \vrf/regTable[3][144] ) );
  LHQD1BWP \vrf/regTable_reg[3][145]  ( .E(n5250), .D(\vrf/N164 ), .Q(
        \vrf/regTable[3][145] ) );
  LHQD1BWP \vrf/regTable_reg[3][146]  ( .E(n5251), .D(\vrf/N165 ), .Q(
        \vrf/regTable[3][146] ) );
  LHQD1BWP \vrf/regTable_reg[3][147]  ( .E(n5251), .D(\vrf/N166 ), .Q(
        \vrf/regTable[3][147] ) );
  LHQD1BWP \vrf/regTable_reg[3][148]  ( .E(n5251), .D(\vrf/N167 ), .Q(
        \vrf/regTable[3][148] ) );
  LHQD1BWP \vrf/regTable_reg[3][149]  ( .E(n5251), .D(\vrf/N168 ), .Q(
        \vrf/regTable[3][149] ) );
  LHQD1BWP \vrf/regTable_reg[3][150]  ( .E(n5251), .D(\vrf/N169 ), .Q(
        \vrf/regTable[3][150] ) );
  LHQD1BWP \vrf/regTable_reg[3][151]  ( .E(n5251), .D(\vrf/N170 ), .Q(
        \vrf/regTable[3][151] ) );
  LHQD1BWP \vrf/regTable_reg[3][152]  ( .E(n5251), .D(\vrf/N171 ), .Q(
        \vrf/regTable[3][152] ) );
  LHQD1BWP \vrf/regTable_reg[3][153]  ( .E(n5251), .D(\vrf/N172 ), .Q(
        \vrf/regTable[3][153] ) );
  LHQD1BWP \vrf/regTable_reg[3][154]  ( .E(n5251), .D(\vrf/N173 ), .Q(
        \vrf/regTable[3][154] ) );
  LHQD1BWP \vrf/regTable_reg[3][155]  ( .E(n5251), .D(\vrf/N174 ), .Q(
        \vrf/regTable[3][155] ) );
  LHQD1BWP \vrf/regTable_reg[3][156]  ( .E(n5251), .D(\vrf/N175 ), .Q(
        \vrf/regTable[3][156] ) );
  LHQD1BWP \vrf/regTable_reg[3][157]  ( .E(n5251), .D(\vrf/N176 ), .Q(
        \vrf/regTable[3][157] ) );
  LHQD1BWP \vrf/regTable_reg[3][158]  ( .E(n5252), .D(\vrf/N177 ), .Q(
        \vrf/regTable[3][158] ) );
  LHQD1BWP \vrf/regTable_reg[3][159]  ( .E(n5252), .D(\vrf/N178 ), .Q(
        \vrf/regTable[3][159] ) );
  LHQD1BWP \vrf/regTable_reg[3][160]  ( .E(n5252), .D(\vrf/N179 ), .Q(
        \vrf/regTable[3][160] ) );
  LHQD1BWP \vrf/regTable_reg[3][161]  ( .E(n5252), .D(\vrf/N180 ), .Q(
        \vrf/regTable[3][161] ) );
  LHQD1BWP \vrf/regTable_reg[3][162]  ( .E(n5252), .D(\vrf/N181 ), .Q(
        \vrf/regTable[3][162] ) );
  LHQD1BWP \vrf/regTable_reg[3][163]  ( .E(n5252), .D(\vrf/N182 ), .Q(
        \vrf/regTable[3][163] ) );
  LHQD1BWP \vrf/regTable_reg[3][164]  ( .E(n5252), .D(\vrf/N183 ), .Q(
        \vrf/regTable[3][164] ) );
  LHQD1BWP \vrf/regTable_reg[3][165]  ( .E(n5252), .D(\vrf/N184 ), .Q(
        \vrf/regTable[3][165] ) );
  LHQD1BWP \vrf/regTable_reg[3][166]  ( .E(n5252), .D(\vrf/N185 ), .Q(
        \vrf/regTable[3][166] ) );
  LHQD1BWP \vrf/regTable_reg[3][167]  ( .E(n5252), .D(\vrf/N186 ), .Q(
        \vrf/regTable[3][167] ) );
  LHQD1BWP \vrf/regTable_reg[3][168]  ( .E(n5252), .D(\vrf/N187 ), .Q(
        \vrf/regTable[3][168] ) );
  LHQD1BWP \vrf/regTable_reg[3][169]  ( .E(n5252), .D(\vrf/N188 ), .Q(
        \vrf/regTable[3][169] ) );
  LHQD1BWP \vrf/regTable_reg[3][170]  ( .E(n5253), .D(\vrf/N189 ), .Q(
        \vrf/regTable[3][170] ) );
  LHQD1BWP \vrf/regTable_reg[3][171]  ( .E(n5253), .D(\vrf/N190 ), .Q(
        \vrf/regTable[3][171] ) );
  LHQD1BWP \vrf/regTable_reg[3][172]  ( .E(n5253), .D(\vrf/N191 ), .Q(
        \vrf/regTable[3][172] ) );
  LHQD1BWP \vrf/regTable_reg[3][173]  ( .E(n5253), .D(\vrf/N192 ), .Q(
        \vrf/regTable[3][173] ) );
  LHQD1BWP \vrf/regTable_reg[3][174]  ( .E(n5253), .D(\vrf/N193 ), .Q(
        \vrf/regTable[3][174] ) );
  LHQD1BWP \vrf/regTable_reg[3][175]  ( .E(n5253), .D(\vrf/N194 ), .Q(
        \vrf/regTable[3][175] ) );
  LHQD1BWP \vrf/regTable_reg[3][176]  ( .E(n5253), .D(\vrf/N195 ), .Q(
        \vrf/regTable[3][176] ) );
  LHQD1BWP \vrf/regTable_reg[3][177]  ( .E(n5253), .D(\vrf/N196 ), .Q(
        \vrf/regTable[3][177] ) );
  LHQD1BWP \vrf/regTable_reg[3][178]  ( .E(n5253), .D(\vrf/N197 ), .Q(
        \vrf/regTable[3][178] ) );
  LHQD1BWP \vrf/regTable_reg[3][179]  ( .E(n5253), .D(\vrf/N198 ), .Q(
        \vrf/regTable[3][179] ) );
  LHQD1BWP \vrf/regTable_reg[3][180]  ( .E(n5253), .D(\vrf/N199 ), .Q(
        \vrf/regTable[3][180] ) );
  LHQD1BWP \vrf/regTable_reg[3][181]  ( .E(n5253), .D(\vrf/N200 ), .Q(
        \vrf/regTable[3][181] ) );
  LHQD1BWP \vrf/regTable_reg[3][182]  ( .E(n5254), .D(\vrf/N201 ), .Q(
        \vrf/regTable[3][182] ) );
  LHQD1BWP \vrf/regTable_reg[3][183]  ( .E(n5254), .D(\vrf/N202 ), .Q(
        \vrf/regTable[3][183] ) );
  LHQD1BWP \vrf/regTable_reg[3][184]  ( .E(n5254), .D(\vrf/N203 ), .Q(
        \vrf/regTable[3][184] ) );
  LHQD1BWP \vrf/regTable_reg[3][185]  ( .E(n5254), .D(\vrf/N204 ), .Q(
        \vrf/regTable[3][185] ) );
  LHQD1BWP \vrf/regTable_reg[3][186]  ( .E(n5254), .D(\vrf/N205 ), .Q(
        \vrf/regTable[3][186] ) );
  LHQD1BWP \vrf/regTable_reg[3][187]  ( .E(n5254), .D(\vrf/N206 ), .Q(
        \vrf/regTable[3][187] ) );
  LHQD1BWP \vrf/regTable_reg[3][188]  ( .E(n5254), .D(\vrf/N207 ), .Q(
        \vrf/regTable[3][188] ) );
  LHQD1BWP \vrf/regTable_reg[3][189]  ( .E(n5254), .D(\vrf/N208 ), .Q(
        \vrf/regTable[3][189] ) );
  LHQD1BWP \vrf/regTable_reg[3][190]  ( .E(n5254), .D(\vrf/N209 ), .Q(
        \vrf/regTable[3][190] ) );
  LHQD1BWP \vrf/regTable_reg[3][191]  ( .E(n5254), .D(\vrf/N210 ), .Q(
        \vrf/regTable[3][191] ) );
  LHQD1BWP \vrf/regTable_reg[3][192]  ( .E(n5254), .D(\vrf/N211 ), .Q(
        \vrf/regTable[3][192] ) );
  LHQD1BWP \vrf/regTable_reg[3][193]  ( .E(n5254), .D(\vrf/N212 ), .Q(
        \vrf/regTable[3][193] ) );
  LHQD1BWP \vrf/regTable_reg[3][194]  ( .E(n5255), .D(\vrf/N213 ), .Q(
        \vrf/regTable[3][194] ) );
  LHQD1BWP \vrf/regTable_reg[3][195]  ( .E(n5255), .D(\vrf/N214 ), .Q(
        \vrf/regTable[3][195] ) );
  LHQD1BWP \vrf/regTable_reg[3][196]  ( .E(n5255), .D(\vrf/N215 ), .Q(
        \vrf/regTable[3][196] ) );
  LHQD1BWP \vrf/regTable_reg[3][197]  ( .E(n5255), .D(\vrf/N216 ), .Q(
        \vrf/regTable[3][197] ) );
  LHQD1BWP \vrf/regTable_reg[3][198]  ( .E(n5255), .D(\vrf/N218 ), .Q(
        \vrf/regTable[3][198] ) );
  LHQD1BWP \vrf/regTable_reg[3][199]  ( .E(n5255), .D(\vrf/N219 ), .Q(
        \vrf/regTable[3][199] ) );
  LHQD1BWP \vrf/regTable_reg[3][200]  ( .E(n5255), .D(\vrf/N220 ), .Q(
        \vrf/regTable[3][200] ) );
  LHQD1BWP \vrf/regTable_reg[3][201]  ( .E(n5255), .D(\vrf/N221 ), .Q(
        \vrf/regTable[3][201] ) );
  LHQD1BWP \vrf/regTable_reg[3][202]  ( .E(n5255), .D(\vrf/N222 ), .Q(
        \vrf/regTable[3][202] ) );
  LHQD1BWP \vrf/regTable_reg[3][203]  ( .E(n5255), .D(\vrf/N223 ), .Q(
        \vrf/regTable[3][203] ) );
  LHQD1BWP \vrf/regTable_reg[3][204]  ( .E(n5255), .D(\vrf/N224 ), .Q(
        \vrf/regTable[3][204] ) );
  LHQD1BWP \vrf/regTable_reg[3][205]  ( .E(n5255), .D(\vrf/N225 ), .Q(
        \vrf/regTable[3][205] ) );
  LHQD1BWP \vrf/regTable_reg[3][206]  ( .E(n5256), .D(\vrf/N226 ), .Q(
        \vrf/regTable[3][206] ) );
  LHQD1BWP \vrf/regTable_reg[3][207]  ( .E(n5256), .D(\vrf/N227 ), .Q(
        \vrf/regTable[3][207] ) );
  LHQD1BWP \vrf/regTable_reg[3][208]  ( .E(n5256), .D(\vrf/N228 ), .Q(
        \vrf/regTable[3][208] ) );
  LHQD1BWP \vrf/regTable_reg[3][209]  ( .E(n5256), .D(\vrf/N229 ), .Q(
        \vrf/regTable[3][209] ) );
  LHQD1BWP \vrf/regTable_reg[3][210]  ( .E(n5256), .D(\vrf/N230 ), .Q(
        \vrf/regTable[3][210] ) );
  LHQD1BWP \vrf/regTable_reg[3][211]  ( .E(n5256), .D(\vrf/N231 ), .Q(
        \vrf/regTable[3][211] ) );
  LHQD1BWP \vrf/regTable_reg[3][212]  ( .E(n5256), .D(\vrf/N232 ), .Q(
        \vrf/regTable[3][212] ) );
  LHQD1BWP \vrf/regTable_reg[3][213]  ( .E(n5256), .D(\vrf/N233 ), .Q(
        \vrf/regTable[3][213] ) );
  LHQD1BWP \vrf/regTable_reg[3][214]  ( .E(n5256), .D(\vrf/N234 ), .Q(
        \vrf/regTable[3][214] ) );
  LHQD1BWP \vrf/regTable_reg[3][215]  ( .E(n5256), .D(\vrf/N235 ), .Q(
        \vrf/regTable[3][215] ) );
  LHQD1BWP \vrf/regTable_reg[3][216]  ( .E(n5256), .D(\vrf/N236 ), .Q(
        \vrf/regTable[3][216] ) );
  LHQD1BWP \vrf/regTable_reg[3][217]  ( .E(n5256), .D(\vrf/N237 ), .Q(
        \vrf/regTable[3][217] ) );
  LHQD1BWP \vrf/regTable_reg[3][218]  ( .E(n5257), .D(\vrf/N238 ), .Q(
        \vrf/regTable[3][218] ) );
  LHQD1BWP \vrf/regTable_reg[3][219]  ( .E(n5257), .D(\vrf/N239 ), .Q(
        \vrf/regTable[3][219] ) );
  LHQD1BWP \vrf/regTable_reg[3][220]  ( .E(n5257), .D(\vrf/N240 ), .Q(
        \vrf/regTable[3][220] ) );
  LHQD1BWP \vrf/regTable_reg[3][221]  ( .E(n5257), .D(\vrf/N241 ), .Q(
        \vrf/regTable[3][221] ) );
  LHQD1BWP \vrf/regTable_reg[3][222]  ( .E(n5257), .D(\vrf/N242 ), .Q(
        \vrf/regTable[3][222] ) );
  LHQD1BWP \vrf/regTable_reg[3][223]  ( .E(n5257), .D(\vrf/N243 ), .Q(
        \vrf/regTable[3][223] ) );
  LHQD1BWP \vrf/regTable_reg[3][224]  ( .E(n5257), .D(\vrf/N244 ), .Q(
        \vrf/regTable[3][224] ) );
  LHQD1BWP \vrf/regTable_reg[3][225]  ( .E(n5257), .D(\vrf/N245 ), .Q(
        \vrf/regTable[3][225] ) );
  LHQD1BWP \vrf/regTable_reg[3][226]  ( .E(n5257), .D(\vrf/N246 ), .Q(
        \vrf/regTable[3][226] ) );
  LHQD1BWP \vrf/regTable_reg[3][227]  ( .E(n5257), .D(\vrf/N247 ), .Q(
        \vrf/regTable[3][227] ) );
  LHQD1BWP \vrf/regTable_reg[3][228]  ( .E(n5257), .D(\vrf/N248 ), .Q(
        \vrf/regTable[3][228] ) );
  LHQD1BWP \vrf/regTable_reg[3][229]  ( .E(n5257), .D(\vrf/N249 ), .Q(
        \vrf/regTable[3][229] ) );
  LHQD1BWP \vrf/regTable_reg[3][230]  ( .E(n5258), .D(\vrf/N250 ), .Q(
        \vrf/regTable[3][230] ) );
  LHQD1BWP \vrf/regTable_reg[3][231]  ( .E(n5258), .D(\vrf/N251 ), .Q(
        \vrf/regTable[3][231] ) );
  LHQD1BWP \vrf/regTable_reg[3][232]  ( .E(n5258), .D(\vrf/N252 ), .Q(
        \vrf/regTable[3][232] ) );
  LHQD1BWP \vrf/regTable_reg[3][233]  ( .E(n5258), .D(\vrf/N253 ), .Q(
        \vrf/regTable[3][233] ) );
  LHQD1BWP \vrf/regTable_reg[3][234]  ( .E(n5258), .D(\vrf/N254 ), .Q(
        \vrf/regTable[3][234] ) );
  LHQD1BWP \vrf/regTable_reg[3][235]  ( .E(n5258), .D(\vrf/N255 ), .Q(
        \vrf/regTable[3][235] ) );
  LHQD1BWP \vrf/regTable_reg[3][236]  ( .E(n5258), .D(\vrf/N256 ), .Q(
        \vrf/regTable[3][236] ) );
  LHQD1BWP \vrf/regTable_reg[3][237]  ( .E(n5258), .D(\vrf/N257 ), .Q(
        \vrf/regTable[3][237] ) );
  LHQD1BWP \vrf/regTable_reg[3][238]  ( .E(n5258), .D(\vrf/N258 ), .Q(
        \vrf/regTable[3][238] ) );
  LHQD1BWP \vrf/regTable_reg[3][239]  ( .E(n5258), .D(\vrf/N259 ), .Q(
        \vrf/regTable[3][239] ) );
  LHQD1BWP \vrf/regTable_reg[3][240]  ( .E(n5258), .D(\vrf/N260 ), .Q(
        \vrf/regTable[3][240] ) );
  LHQD1BWP \vrf/regTable_reg[3][241]  ( .E(n5258), .D(\vrf/N261 ), .Q(
        \vrf/regTable[3][241] ) );
  LHQD1BWP \vrf/regTable_reg[3][242]  ( .E(n5259), .D(\vrf/N262 ), .Q(
        \vrf/regTable[3][242] ) );
  LHQD1BWP \vrf/regTable_reg[3][243]  ( .E(n5259), .D(\vrf/N263 ), .Q(
        \vrf/regTable[3][243] ) );
  LHQD1BWP \vrf/regTable_reg[3][244]  ( .E(n5259), .D(\vrf/N264 ), .Q(
        \vrf/regTable[3][244] ) );
  LHQD1BWP \vrf/regTable_reg[3][245]  ( .E(n5259), .D(\vrf/N265 ), .Q(
        \vrf/regTable[3][245] ) );
  LHQD1BWP \vrf/regTable_reg[3][246]  ( .E(n5259), .D(\vrf/N266 ), .Q(
        \vrf/regTable[3][246] ) );
  LHQD1BWP \vrf/regTable_reg[3][247]  ( .E(n5259), .D(\vrf/N267 ), .Q(
        \vrf/regTable[3][247] ) );
  LHQD1BWP \vrf/regTable_reg[3][248]  ( .E(n5259), .D(\vrf/N268 ), .Q(
        \vrf/regTable[3][248] ) );
  LHQD1BWP \vrf/regTable_reg[3][249]  ( .E(n5259), .D(\vrf/N269 ), .Q(
        \vrf/regTable[3][249] ) );
  LHQD1BWP \vrf/regTable_reg[3][250]  ( .E(n5259), .D(\vrf/N270 ), .Q(
        \vrf/regTable[3][250] ) );
  LHQD1BWP \vrf/regTable_reg[3][251]  ( .E(n5259), .D(\vrf/N271 ), .Q(
        \vrf/regTable[3][251] ) );
  LHQD1BWP \vrf/regTable_reg[3][252]  ( .E(n5259), .D(\vrf/N272 ), .Q(
        \vrf/regTable[3][252] ) );
  LHQD1BWP \vrf/regTable_reg[3][253]  ( .E(n5259), .D(\vrf/N273 ), .Q(
        \vrf/regTable[3][253] ) );
  LHQD1BWP \wrAddr_reg[0]  ( .E(N4366), .D(addrDst[0]), .Q(\srf/N15 ) );
  LHQD1BWP \op1_reg[11]  ( .E(N4102), .D(N4081), .Q(op1[11]) );
  LHQD1BWP \op2_reg[12]  ( .E(N4102), .D(N4098), .Q(op2[12]) );
  LNQD1BWP \scalarToLoad_reg[10]  ( .D(N1757), .EN(n2522), .Q(scalarToLoad[10]) );
  LNQD1BWP \instrIn_reg[15]  ( .D(DataIn[15]), .EN(n3262), .Q(code[3]) );
  LHQD1BWP \op2_reg[11]  ( .E(N4102), .D(N4097), .Q(op2[11]) );
  LHQD1BWP \op1_reg[10]  ( .E(N4102), .D(N4080), .Q(op1[10]) );
  LHQD1BWP \op1_reg[12]  ( .E(N4102), .D(N4082), .Q(op1[12]) );
  LHQD1BWP \op1_reg[15]  ( .E(N4102), .D(N4085), .Q(op1[15]) );
  LHQD1BWP \srf/regTable_reg[6][0]  ( .E(\srf/N53 ), .D(\srf/N37 ), .Q(
        \srf/regTable[6][0] ) );
  LHQD1BWP \srf/regTable_reg[6][1]  ( .E(\srf/N53 ), .D(\srf/N38 ), .Q(
        \srf/regTable[6][1] ) );
  LHQD1BWP \srf/regTable_reg[6][2]  ( .E(\srf/N53 ), .D(\srf/N39 ), .Q(
        \srf/regTable[6][2] ) );
  LHQD1BWP \srf/regTable_reg[6][3]  ( .E(\srf/N53 ), .D(\srf/N40 ), .Q(
        \srf/regTable[6][3] ) );
  LHQD1BWP \srf/regTable_reg[6][4]  ( .E(\srf/N53 ), .D(\srf/N41 ), .Q(
        \srf/regTable[6][4] ) );
  LHQD1BWP \srf/regTable_reg[6][5]  ( .E(\srf/N53 ), .D(\srf/N42 ), .Q(
        \srf/regTable[6][5] ) );
  LHQD1BWP \srf/regTable_reg[6][6]  ( .E(\srf/N53 ), .D(\srf/N43 ), .Q(
        \srf/regTable[6][6] ) );
  LHQD1BWP \srf/regTable_reg[6][7]  ( .E(\srf/N53 ), .D(\srf/N44 ), .Q(
        \srf/regTable[6][7] ) );
  LHQD1BWP \srf/regTable_reg[6][8]  ( .E(\srf/N53 ), .D(\srf/N45 ), .Q(
        \srf/regTable[6][8] ) );
  LHQD1BWP \srf/regTable_reg[6][9]  ( .E(\srf/N53 ), .D(\srf/N46 ), .Q(
        \srf/regTable[6][9] ) );
  LHQD1BWP \srf/regTable_reg[6][10]  ( .E(\srf/N53 ), .D(\srf/N47 ), .Q(
        \srf/regTable[6][10] ) );
  LHQD1BWP \srf/regTable_reg[6][11]  ( .E(\srf/N53 ), .D(\srf/N48 ), .Q(
        \srf/regTable[6][11] ) );
  LHQD1BWP \srf/regTable_reg[6][12]  ( .E(\srf/N53 ), .D(\srf/N49 ), .Q(
        \srf/regTable[6][12] ) );
  LHQD1BWP \srf/regTable_reg[6][13]  ( .E(\srf/N53 ), .D(\srf/N50 ), .Q(
        \srf/regTable[6][13] ) );
  LHQD1BWP \srf/regTable_reg[6][14]  ( .E(\srf/N53 ), .D(\srf/N51 ), .Q(
        \srf/regTable[6][14] ) );
  LHQD1BWP \srf/regTable_reg[6][15]  ( .E(\srf/N53 ), .D(\srf/N52 ), .Q(
        \srf/regTable[6][15] ) );
  LHQD1BWP \srf/regTable_reg[4][0]  ( .E(\srf/N55 ), .D(\srf/N37 ), .Q(
        \srf/regTable[4][0] ) );
  LHQD1BWP \srf/regTable_reg[4][1]  ( .E(\srf/N55 ), .D(\srf/N38 ), .Q(
        \srf/regTable[4][1] ) );
  LHQD1BWP \srf/regTable_reg[4][2]  ( .E(\srf/N55 ), .D(\srf/N39 ), .Q(
        \srf/regTable[4][2] ) );
  LHQD1BWP \srf/regTable_reg[4][3]  ( .E(\srf/N55 ), .D(\srf/N40 ), .Q(
        \srf/regTable[4][3] ) );
  LHQD1BWP \srf/regTable_reg[4][4]  ( .E(\srf/N55 ), .D(\srf/N41 ), .Q(
        \srf/regTable[4][4] ) );
  LHQD1BWP \srf/regTable_reg[4][5]  ( .E(\srf/N55 ), .D(\srf/N42 ), .Q(
        \srf/regTable[4][5] ) );
  LHQD1BWP \srf/regTable_reg[4][6]  ( .E(\srf/N55 ), .D(\srf/N43 ), .Q(
        \srf/regTable[4][6] ) );
  LHQD1BWP \srf/regTable_reg[4][7]  ( .E(\srf/N55 ), .D(\srf/N44 ), .Q(
        \srf/regTable[4][7] ) );
  LHQD1BWP \srf/regTable_reg[4][8]  ( .E(\srf/N55 ), .D(\srf/N45 ), .Q(
        \srf/regTable[4][8] ) );
  LHQD1BWP \srf/regTable_reg[4][9]  ( .E(\srf/N55 ), .D(\srf/N46 ), .Q(
        \srf/regTable[4][9] ) );
  LHQD1BWP \srf/regTable_reg[4][10]  ( .E(\srf/N55 ), .D(\srf/N47 ), .Q(
        \srf/regTable[4][10] ) );
  LHQD1BWP \srf/regTable_reg[4][11]  ( .E(\srf/N55 ), .D(\srf/N48 ), .Q(
        \srf/regTable[4][11] ) );
  LHQD1BWP \srf/regTable_reg[4][12]  ( .E(\srf/N55 ), .D(\srf/N49 ), .Q(
        \srf/regTable[4][12] ) );
  LHQD1BWP \srf/regTable_reg[4][13]  ( .E(\srf/N55 ), .D(\srf/N50 ), .Q(
        \srf/regTable[4][13] ) );
  LHQD1BWP \srf/regTable_reg[4][14]  ( .E(\srf/N55 ), .D(\srf/N51 ), .Q(
        \srf/regTable[4][14] ) );
  LHQD1BWP \srf/regTable_reg[4][15]  ( .E(\srf/N55 ), .D(\srf/N52 ), .Q(
        \srf/regTable[4][15] ) );
  LHQD1BWP \srf/regTable_reg[2][0]  ( .E(\srf/N57 ), .D(\srf/N37 ), .Q(
        \srf/regTable[2][0] ) );
  LHQD1BWP \srf/regTable_reg[2][1]  ( .E(\srf/N57 ), .D(\srf/N38 ), .Q(
        \srf/regTable[2][1] ) );
  LHQD1BWP \srf/regTable_reg[2][2]  ( .E(\srf/N57 ), .D(\srf/N39 ), .Q(
        \srf/regTable[2][2] ) );
  LHQD1BWP \srf/regTable_reg[2][3]  ( .E(\srf/N57 ), .D(\srf/N40 ), .Q(
        \srf/regTable[2][3] ) );
  LHQD1BWP \srf/regTable_reg[2][4]  ( .E(\srf/N57 ), .D(\srf/N41 ), .Q(
        \srf/regTable[2][4] ) );
  LHQD1BWP \srf/regTable_reg[2][5]  ( .E(\srf/N57 ), .D(\srf/N42 ), .Q(
        \srf/regTable[2][5] ) );
  LHQD1BWP \srf/regTable_reg[2][6]  ( .E(\srf/N57 ), .D(\srf/N43 ), .Q(
        \srf/regTable[2][6] ) );
  LHQD1BWP \srf/regTable_reg[2][7]  ( .E(\srf/N57 ), .D(\srf/N44 ), .Q(
        \srf/regTable[2][7] ) );
  LHQD1BWP \srf/regTable_reg[2][8]  ( .E(\srf/N57 ), .D(\srf/N45 ), .Q(
        \srf/regTable[2][8] ) );
  LHQD1BWP \srf/regTable_reg[2][9]  ( .E(\srf/N57 ), .D(\srf/N46 ), .Q(
        \srf/regTable[2][9] ) );
  LHQD1BWP \srf/regTable_reg[2][10]  ( .E(\srf/N57 ), .D(\srf/N47 ), .Q(
        \srf/regTable[2][10] ) );
  LHQD1BWP \srf/regTable_reg[2][11]  ( .E(\srf/N57 ), .D(\srf/N48 ), .Q(
        \srf/regTable[2][11] ) );
  LHQD1BWP \srf/regTable_reg[2][12]  ( .E(\srf/N57 ), .D(\srf/N49 ), .Q(
        \srf/regTable[2][12] ) );
  LHQD1BWP \srf/regTable_reg[2][13]  ( .E(\srf/N57 ), .D(\srf/N50 ), .Q(
        \srf/regTable[2][13] ) );
  LHQD1BWP \srf/regTable_reg[2][14]  ( .E(\srf/N57 ), .D(\srf/N51 ), .Q(
        \srf/regTable[2][14] ) );
  LHQD1BWP \srf/regTable_reg[2][15]  ( .E(\srf/N57 ), .D(\srf/N52 ), .Q(
        \srf/regTable[2][15] ) );
  LHQD1BWP \srf/regTable_reg[0][0]  ( .E(\srf/N59 ), .D(\srf/N37 ), .Q(
        \srf/regTable[0][0] ) );
  LHQD1BWP \srf/regTable_reg[0][1]  ( .E(\srf/N59 ), .D(\srf/N38 ), .Q(
        \srf/regTable[0][1] ) );
  LHQD1BWP \srf/regTable_reg[0][2]  ( .E(\srf/N59 ), .D(\srf/N39 ), .Q(
        \srf/regTable[0][2] ) );
  LHQD1BWP \srf/regTable_reg[0][3]  ( .E(\srf/N59 ), .D(\srf/N40 ), .Q(
        \srf/regTable[0][3] ) );
  LHQD1BWP \srf/regTable_reg[0][4]  ( .E(\srf/N59 ), .D(\srf/N41 ), .Q(
        \srf/regTable[0][4] ) );
  LHQD1BWP \srf/regTable_reg[0][5]  ( .E(\srf/N59 ), .D(\srf/N42 ), .Q(
        \srf/regTable[0][5] ) );
  LHQD1BWP \srf/regTable_reg[0][6]  ( .E(\srf/N59 ), .D(\srf/N43 ), .Q(
        \srf/regTable[0][6] ) );
  LHQD1BWP \srf/regTable_reg[0][7]  ( .E(\srf/N59 ), .D(\srf/N44 ), .Q(
        \srf/regTable[0][7] ) );
  LHQD1BWP \srf/regTable_reg[0][8]  ( .E(\srf/N59 ), .D(\srf/N45 ), .Q(
        \srf/regTable[0][8] ) );
  LHQD1BWP \srf/regTable_reg[0][9]  ( .E(\srf/N59 ), .D(\srf/N46 ), .Q(
        \srf/regTable[0][9] ) );
  LHQD1BWP \srf/regTable_reg[0][10]  ( .E(\srf/N59 ), .D(\srf/N47 ), .Q(
        \srf/regTable[0][10] ) );
  LHQD1BWP \srf/regTable_reg[0][11]  ( .E(\srf/N59 ), .D(\srf/N48 ), .Q(
        \srf/regTable[0][11] ) );
  LHQD1BWP \srf/regTable_reg[0][12]  ( .E(\srf/N59 ), .D(\srf/N49 ), .Q(
        \srf/regTable[0][12] ) );
  LHQD1BWP \srf/regTable_reg[0][13]  ( .E(\srf/N59 ), .D(\srf/N50 ), .Q(
        \srf/regTable[0][13] ) );
  LHQD1BWP \srf/regTable_reg[0][14]  ( .E(\srf/N59 ), .D(\srf/N51 ), .Q(
        \srf/regTable[0][14] ) );
  LHQD1BWP \srf/regTable_reg[0][15]  ( .E(\srf/N59 ), .D(\srf/N52 ), .Q(
        \srf/regTable[0][15] ) );
  LNQD1BWP \instrIn_reg[13]  ( .D(DataIn[13]), .EN(n3262), .Q(code[1]) );
  LHQD1BWP \op1_reg[13]  ( .E(N4102), .D(N4083), .Q(op1[13]) );
  LHQD1BWP \srf/regTable_reg[5][0]  ( .E(\srf/N54 ), .D(\srf/N37 ), .Q(
        \srf/regTable[5][0] ) );
  LHQD1BWP \srf/regTable_reg[5][1]  ( .E(\srf/N54 ), .D(\srf/N38 ), .Q(
        \srf/regTable[5][1] ) );
  LHQD1BWP \srf/regTable_reg[5][2]  ( .E(\srf/N54 ), .D(\srf/N39 ), .Q(
        \srf/regTable[5][2] ) );
  LHQD1BWP \srf/regTable_reg[5][3]  ( .E(\srf/N54 ), .D(\srf/N40 ), .Q(
        \srf/regTable[5][3] ) );
  LHQD1BWP \srf/regTable_reg[5][4]  ( .E(\srf/N54 ), .D(\srf/N41 ), .Q(
        \srf/regTable[5][4] ) );
  LHQD1BWP \srf/regTable_reg[5][5]  ( .E(\srf/N54 ), .D(\srf/N42 ), .Q(
        \srf/regTable[5][5] ) );
  LHQD1BWP \srf/regTable_reg[5][6]  ( .E(\srf/N54 ), .D(\srf/N43 ), .Q(
        \srf/regTable[5][6] ) );
  LHQD1BWP \srf/regTable_reg[5][7]  ( .E(\srf/N54 ), .D(\srf/N44 ), .Q(
        \srf/regTable[5][7] ) );
  LHQD1BWP \srf/regTable_reg[5][8]  ( .E(\srf/N54 ), .D(\srf/N45 ), .Q(
        \srf/regTable[5][8] ) );
  LHQD1BWP \srf/regTable_reg[5][9]  ( .E(\srf/N54 ), .D(\srf/N46 ), .Q(
        \srf/regTable[5][9] ) );
  LHQD1BWP \srf/regTable_reg[1][0]  ( .E(\srf/N58 ), .D(\srf/N37 ), .Q(
        \srf/regTable[1][0] ) );
  LHQD1BWP \srf/regTable_reg[1][1]  ( .E(\srf/N58 ), .D(\srf/N38 ), .Q(
        \srf/regTable[1][1] ) );
  LHQD1BWP \srf/regTable_reg[1][2]  ( .E(\srf/N58 ), .D(\srf/N39 ), .Q(
        \srf/regTable[1][2] ) );
  LHQD1BWP \srf/regTable_reg[1][3]  ( .E(\srf/N58 ), .D(\srf/N40 ), .Q(
        \srf/regTable[1][3] ) );
  LHQD1BWP \srf/regTable_reg[1][4]  ( .E(\srf/N58 ), .D(\srf/N41 ), .Q(
        \srf/regTable[1][4] ) );
  LHQD1BWP \srf/regTable_reg[1][5]  ( .E(\srf/N58 ), .D(\srf/N42 ), .Q(
        \srf/regTable[1][5] ) );
  LHQD1BWP \srf/regTable_reg[1][6]  ( .E(\srf/N58 ), .D(\srf/N43 ), .Q(
        \srf/regTable[1][6] ) );
  LHQD1BWP \srf/regTable_reg[1][7]  ( .E(\srf/N58 ), .D(\srf/N44 ), .Q(
        \srf/regTable[1][7] ) );
  LHQD1BWP \srf/regTable_reg[1][8]  ( .E(\srf/N58 ), .D(\srf/N45 ), .Q(
        \srf/regTable[1][8] ) );
  LHQD1BWP \srf/regTable_reg[1][9]  ( .E(\srf/N58 ), .D(\srf/N46 ), .Q(
        \srf/regTable[1][9] ) );
  LNQD1BWP \scalarToLoad_reg[12]  ( .D(N1759), .EN(n2522), .Q(scalarToLoad[12]) );
  LHQD1BWP \op2_reg[10]  ( .E(N4102), .D(N4096), .Q(op2[10]) );
  LHQD1BWP \srf/regTable_reg[7][0]  ( .E(\srf/N36 ), .D(\srf/N37 ), .Q(
        \srf/regTable[7][0] ) );
  LHQD1BWP \srf/regTable_reg[7][1]  ( .E(\srf/N36 ), .D(\srf/N38 ), .Q(
        \srf/regTable[7][1] ) );
  LHQD1BWP \srf/regTable_reg[7][2]  ( .E(\srf/N36 ), .D(\srf/N39 ), .Q(
        \srf/regTable[7][2] ) );
  LHQD1BWP \srf/regTable_reg[7][3]  ( .E(\srf/N36 ), .D(\srf/N40 ), .Q(
        \srf/regTable[7][3] ) );
  LHQD1BWP \srf/regTable_reg[7][4]  ( .E(\srf/N36 ), .D(\srf/N41 ), .Q(
        \srf/regTable[7][4] ) );
  LHQD1BWP \srf/regTable_reg[7][5]  ( .E(\srf/N36 ), .D(\srf/N42 ), .Q(
        \srf/regTable[7][5] ) );
  LHQD1BWP \srf/regTable_reg[7][6]  ( .E(\srf/N36 ), .D(\srf/N43 ), .Q(
        \srf/regTable[7][6] ) );
  LHQD1BWP \srf/regTable_reg[7][7]  ( .E(\srf/N36 ), .D(\srf/N44 ), .Q(
        \srf/regTable[7][7] ) );
  LHQD1BWP \srf/regTable_reg[7][8]  ( .E(\srf/N36 ), .D(\srf/N45 ), .Q(
        \srf/regTable[7][8] ) );
  LHQD1BWP \srf/regTable_reg[7][9]  ( .E(\srf/N36 ), .D(\srf/N46 ), .Q(
        \srf/regTable[7][9] ) );
  LHQD1BWP \srf/regTable_reg[3][0]  ( .E(\srf/N56 ), .D(\srf/N37 ), .Q(
        \srf/regTable[3][0] ) );
  LHQD1BWP \srf/regTable_reg[3][1]  ( .E(\srf/N56 ), .D(\srf/N38 ), .Q(
        \srf/regTable[3][1] ) );
  LHQD1BWP \srf/regTable_reg[3][2]  ( .E(\srf/N56 ), .D(\srf/N39 ), .Q(
        \srf/regTable[3][2] ) );
  LHQD1BWP \srf/regTable_reg[3][3]  ( .E(\srf/N56 ), .D(\srf/N40 ), .Q(
        \srf/regTable[3][3] ) );
  LHQD1BWP \srf/regTable_reg[3][4]  ( .E(\srf/N56 ), .D(\srf/N41 ), .Q(
        \srf/regTable[3][4] ) );
  LHQD1BWP \srf/regTable_reg[3][5]  ( .E(\srf/N56 ), .D(\srf/N42 ), .Q(
        \srf/regTable[3][5] ) );
  LHQD1BWP \srf/regTable_reg[3][6]  ( .E(\srf/N56 ), .D(\srf/N43 ), .Q(
        \srf/regTable[3][6] ) );
  LHQD1BWP \srf/regTable_reg[3][7]  ( .E(\srf/N56 ), .D(\srf/N44 ), .Q(
        \srf/regTable[3][7] ) );
  LHQD1BWP \srf/regTable_reg[3][8]  ( .E(\srf/N56 ), .D(\srf/N45 ), .Q(
        \srf/regTable[3][8] ) );
  LHQD1BWP \srf/regTable_reg[3][9]  ( .E(\srf/N56 ), .D(\srf/N46 ), .Q(
        \srf/regTable[3][9] ) );
  LHQD1BWP \op2_reg[13]  ( .E(N4102), .D(N4099), .Q(op2[13]) );
  LNQD1BWP \instrIn_reg[12]  ( .D(DataIn[12]), .EN(n3262), .Q(code[0]) );
  LNQD1BWP \scalarToLoad_reg[13]  ( .D(N1760), .EN(n2522), .Q(scalarToLoad[13]) );
  LNQD1BWP \scalarToLoad_reg[14]  ( .D(N1761), .EN(n2522), .Q(scalarToLoad[14]) );
  LNQD1BWP \instrIn_reg[14]  ( .D(DataIn[14]), .EN(n3262), .Q(code[2]) );
  LHQD1BWP \op1_reg[14]  ( .E(N4102), .D(N4084), .Q(\alu/N851 ) );
  LND1BWP \scalarToLoad_reg[9]  ( .D(N1756), .EN(n2522), .Q(scalarToLoad[9]), 
        .QN(n3390) );
  LND1BWP \scalarToLoad_reg[8]  ( .D(N1755), .EN(n2522), .Q(scalarToLoad[8]), 
        .QN(n3391) );
  LND1BWP \scalarToLoad_reg[0]  ( .D(N1747), .EN(n2522), .Q(scalarToLoad[0]), 
        .QN(n3389) );
  LND1BWP \scalarToLoad_reg[2]  ( .D(N1749), .EN(n2522), .Q(scalarToLoad[2]), 
        .QN(n3387) );
  LND1BWP \scalarToLoad_reg[1]  ( .D(N1748), .EN(n2522), .Q(scalarToLoad[1]), 
        .QN(n3388) );
  LHQD1BWP \func_reg[1]  ( .E(n3368), .D(code[1]), .Q(func[1]) );
  LND1BWP \scalarToLoad_reg[7]  ( .D(N1754), .EN(n2522), .Q(scalarToLoad[7]), 
        .QN(n3382) );
  LND1BWP \scalarToLoad_reg[6]  ( .D(N1753), .EN(n2522), .Q(scalarToLoad[6]), 
        .QN(n3383) );
  LND1BWP \scalarToLoad_reg[5]  ( .D(N1752), .EN(n2522), .Q(scalarToLoad[5]), 
        .QN(n3384) );
  LND1BWP \scalarToLoad_reg[4]  ( .D(N1751), .EN(n2522), .Q(scalarToLoad[4]), 
        .QN(n3385) );
  LND1BWP \scalarToLoad_reg[3]  ( .D(N1750), .EN(n2522), .Q(scalarToLoad[3]), 
        .QN(n3386) );
  LHQD1BWP \op2_reg[9]  ( .E(N4102), .D(N4095), .Q(op2[9]) );
  LHQD1BWP \op2_reg[8]  ( .E(N4102), .D(N4094), .Q(op2[8]) );
  LHQD1BWP \op1_reg[9]  ( .E(N4102), .D(N4079), .Q(op1[9]) );
  LHQD1BWP \op1_reg[8]  ( .E(N4102), .D(N4078), .Q(op1[8]) );
  LHD1BWP \op1_reg[7]  ( .E(N4102), .D(N4077), .Q(op1[7]), .QN(n3370) );
  LHQD1BWP \op1_reg[1]  ( .E(N4102), .D(N4071), .Q(op1[1]) );
  LHD1BWP \op1_reg[2]  ( .E(N4102), .D(N4072), .Q(op1[2]), .QN(n3371) );
  LHQD1BWP \op2_reg[1]  ( .E(N4102), .D(N4087), .Q(op2[1]) );
  LHD1BWP \op2_reg[2]  ( .E(N4102), .D(N4088), .Q(op2[2]), .QN(n3379) );
  LHQD1BWP \op2_reg[0]  ( .E(N4102), .D(N4086), .Q(op2[0]) );
  LHD1BWP \op1_reg[6]  ( .E(N4102), .D(N4076), .Q(op1[6]), .QN(n3380) );
  LHD1BWP \op1_reg[4]  ( .E(N4102), .D(N4074), .Q(op1[4]), .QN(n3376) );
  LHD1BWP \op1_reg[3]  ( .E(N4102), .D(N4073), .Q(op1[3]), .QN(n3381) );
  LHD1BWP \op1_reg[5]  ( .E(N4102), .D(N4075), .Q(op1[5]), .QN(n3377) );
  LHD1BWP \op2_reg[6]  ( .E(N4102), .D(N4092), .Q(op2[6]), .QN(n3372) );
  LHD1BWP \op2_reg[5]  ( .E(N4102), .D(N4091), .Q(op2[5]), .QN(n3378) );
  LHD1BWP \op2_reg[4]  ( .E(N4102), .D(N4090), .Q(op2[4]), .QN(n3373) );
  LHD1BWP \op2_reg[3]  ( .E(N4102), .D(N4089), .Q(op2[3]), .QN(n3375) );
  LHD1BWP \op2_reg[7]  ( .E(N4102), .D(N4093), .Q(op2[7]), .QN(n3374) );
  LHQD2BWP \wrAddr_reg[1]  ( .E(N4366), .D(addrDst[1]), .Q(\srf/N16 ) );
  LHQD2BWP \func_reg[2]  ( .E(n3368), .D(code[2]), .Q(func[2]) );
  LHQD2BWP \func_reg[0]  ( .E(n3368), .D(code[0]), .Q(func[0]) );
  LNCNQD1BWP flow_reg ( .D(overflow), .EN(n3266), .CDN(n7436), .Q(V) );
  LHQD1BWP \op1_reg[0]  ( .E(N4102), .D(N4070), .Q(op1[0]) );
  LHQD1BWP overflow_reg ( .E(N4103), .D(N4104), .Q(overflow) );
  LHQD2BWP \func_reg[3]  ( .E(n3368), .D(code[3]), .Q(func[3]) );
  LHQD1BWP \srf/regTable_reg[7][10]  ( .E(\srf/N36 ), .D(\srf/N47 ), .Q(
        \srf/regTable[7][10] ) );
  LHQD1BWP \srf/regTable_reg[7][11]  ( .E(\srf/N36 ), .D(\srf/N48 ), .Q(
        \srf/regTable[7][11] ) );
  LHQD1BWP \srf/regTable_reg[7][12]  ( .E(\srf/N36 ), .D(\srf/N49 ), .Q(
        \srf/regTable[7][12] ) );
  LHQD1BWP \srf/regTable_reg[7][13]  ( .E(\srf/N36 ), .D(\srf/N50 ), .Q(
        \srf/regTable[7][13] ) );
  LHQD1BWP \srf/regTable_reg[7][14]  ( .E(\srf/N36 ), .D(\srf/N51 ), .Q(
        \srf/regTable[7][14] ) );
  LHQD1BWP \srf/regTable_reg[7][15]  ( .E(\srf/N36 ), .D(\srf/N52 ), .Q(
        \srf/regTable[7][15] ) );
  LHQD1BWP \srf/regTable_reg[5][10]  ( .E(\srf/N54 ), .D(\srf/N47 ), .Q(
        \srf/regTable[5][10] ) );
  LHQD1BWP \srf/regTable_reg[5][11]  ( .E(\srf/N54 ), .D(\srf/N48 ), .Q(
        \srf/regTable[5][11] ) );
  LHQD1BWP \srf/regTable_reg[5][12]  ( .E(\srf/N54 ), .D(\srf/N49 ), .Q(
        \srf/regTable[5][12] ) );
  LHQD1BWP \srf/regTable_reg[5][13]  ( .E(\srf/N54 ), .D(\srf/N50 ), .Q(
        \srf/regTable[5][13] ) );
  LHQD1BWP \srf/regTable_reg[5][14]  ( .E(\srf/N54 ), .D(\srf/N51 ), .Q(
        \srf/regTable[5][14] ) );
  LHQD1BWP \srf/regTable_reg[5][15]  ( .E(\srf/N54 ), .D(\srf/N52 ), .Q(
        \srf/regTable[5][15] ) );
  LHQD1BWP \srf/regTable_reg[3][10]  ( .E(\srf/N56 ), .D(\srf/N47 ), .Q(
        \srf/regTable[3][10] ) );
  LHQD1BWP \srf/regTable_reg[3][11]  ( .E(\srf/N56 ), .D(\srf/N48 ), .Q(
        \srf/regTable[3][11] ) );
  LHQD1BWP \srf/regTable_reg[3][12]  ( .E(\srf/N56 ), .D(\srf/N49 ), .Q(
        \srf/regTable[3][12] ) );
  LHQD1BWP \srf/regTable_reg[3][13]  ( .E(\srf/N56 ), .D(\srf/N50 ), .Q(
        \srf/regTable[3][13] ) );
  LHQD1BWP \srf/regTable_reg[3][14]  ( .E(\srf/N56 ), .D(\srf/N51 ), .Q(
        \srf/regTable[3][14] ) );
  LHQD1BWP \srf/regTable_reg[3][15]  ( .E(\srf/N56 ), .D(\srf/N52 ), .Q(
        \srf/regTable[3][15] ) );
  LHQD1BWP \srf/regTable_reg[1][10]  ( .E(\srf/N58 ), .D(\srf/N47 ), .Q(
        \srf/regTable[1][10] ) );
  LHQD1BWP \srf/regTable_reg[1][11]  ( .E(\srf/N58 ), .D(\srf/N48 ), .Q(
        \srf/regTable[1][11] ) );
  LHQD1BWP \srf/regTable_reg[1][12]  ( .E(\srf/N58 ), .D(\srf/N49 ), .Q(
        \srf/regTable[1][12] ) );
  LHQD1BWP \srf/regTable_reg[1][13]  ( .E(\srf/N58 ), .D(\srf/N50 ), .Q(
        \srf/regTable[1][13] ) );
  LHQD1BWP \srf/regTable_reg[1][14]  ( .E(\srf/N58 ), .D(\srf/N51 ), .Q(
        \srf/regTable[1][14] ) );
  LHQD1BWP \srf/regTable_reg[1][15]  ( .E(\srf/N58 ), .D(\srf/N52 ), .Q(
        \srf/regTable[1][15] ) );
  INR3D1BWP U4229 ( .A1(n6052), .B1(n7460), .B2(n6051), .ZN(\alu/N579 ) );
  INR3D1BWP U4230 ( .A1(n6107), .B1(n6104), .B2(\alu/N337 ), .ZN(\alu/N385 )
         );
  INR3D1BWP U4231 ( .A1(n6177), .B1(n7148), .B2(N1418), .ZN(N1466) );
  NR2XD1BWP U4232 ( .A1(n7041), .A2(WR), .ZN(n6171) );
  NR4D1BWP U4233 ( .A1(n7449), .A2(n7448), .A3(N1610), .A4(n7100), .ZN(N1660)
         );
  CKND2BWP U4234 ( .I(n5988), .ZN(n5987) );
  CKND2BWP U4235 ( .I(n6023), .ZN(n5947) );
  OAI22D1BWP U4236 ( .A1(n6108), .A2(n6109), .B1(n6110), .B2(n6005), .ZN(n6023) );
  NR3D1BWP U4237 ( .A1(n5929), .A2(n5935), .A3(n5936), .ZN(n5948) );
  AOI22D2BWP U4238 ( .A1(n7074), .A2(n7112), .B1(cycles[0]), .B2(n6215), .ZN(
        N1561) );
  OAI21D1BWP U4239 ( .A1(n7101), .A2(N1610), .B(n6149), .ZN(N1681) );
  INVD1BWP U4240 ( .I(n6172), .ZN(n7456) );
  CKAN2D0BWP U4241 ( .A1(\alu/N477 ), .A2(n5948), .Z(n5912) );
  MUX2D0BWP U4242 ( .I0(n7468), .I1(\alu/N465 ), .S(n5948), .Z(\alu/N520 ) );
  OAI21D1BWP U4243 ( .A1(n6060), .A2(\alu/N529 ), .B(n6053), .ZN(\alu/N600 )
         );
  MUX2D0BWP U4244 ( .I0(\alu/N449 ), .I1(\alu/N469 ), .S(n5948), .Z(n7463) );
  MUX2D0BWP U4245 ( .I0(\alu/N450 ), .I1(\alu/N470 ), .S(n5948), .Z(n7464) );
  MUX2D0BWP U4246 ( .I0(\alu/N454 ), .I1(\alu/N474 ), .S(n5948), .Z(\alu/N529 ) );
  MUX2D0BWP U4247 ( .I0(\alu/N453 ), .I1(\alu/N473 ), .S(n5948), .Z(n7467) );
  CKAN2D1BWP U4248 ( .A1(n6171), .A2(n6205), .Z(n7008) );
  MUX2D0BWP U4249 ( .I0(n7469), .I1(\alu/N464 ), .S(n5948), .Z(\alu/N519 ) );
  OAI21D1BWP U4250 ( .A1(N1417), .A2(n7158), .B(n6174), .ZN(N1487) );
  OAI21D1BWP U4251 ( .A1(\alu/N336 ), .A2(n6140), .B(n6136), .ZN(\alu/N406 )
         );
  IND2D1BWP U4252 ( .A1(N4104), .B1(n6250), .ZN(N4102) );
  MUX2D0BWP U4253 ( .I0(\alu/N447 ), .I1(\alu/N467 ), .S(n5948), .Z(n7461) );
  XOR3D1BWP U4254 ( .A1(n6204), .A2(n7111), .A3(n7110), .Z(N1563) );
  XNR3D1BWP U4255 ( .A1(n6204), .A2(n7118), .A3(N1561), .ZN(N1562) );
  OAI21D1BWP U4256 ( .A1(n7437), .A2(n5530), .B(n7436), .ZN(\srf/N58 ) );
  OAI21D1BWP U4257 ( .A1(n7437), .A2(n5532), .B(n7436), .ZN(\srf/N56 ) );
  OAI21D1BWP U4258 ( .A1(n7437), .A2(n5533), .B(n7436), .ZN(\srf/N54 ) );
  OAI21D1BWP U4259 ( .A1(n7437), .A2(n5534), .B(n7436), .ZN(\srf/N36 ) );
  MUX2D0BWP U4260 ( .I0(\alu/N107 ), .I1(\alu/N216 ), .S(n5947), .Z(
        \U3/U26/Z_15 ) );
  MUX2D0BWP U4261 ( .I0(N1188), .I1(N1297), .S(n5987), .Z(\U3/U7/Z_15 ) );
  MUX2D0BWP U4262 ( .I0(\alu/N106 ), .I1(\alu/N215 ), .S(n5947), .Z(
        \U3/U26/Z_14 ) );
  MUX2D0BWP U4263 ( .I0(N1187), .I1(N1296), .S(n5987), .Z(\U3/U7/Z_14 ) );
  MUX2D0BWP U4264 ( .I0(\alu/N101 ), .I1(\alu/N210 ), .S(n5947), .Z(
        \U3/U26/Z_9 ) );
  MUX2D0BWP U4265 ( .I0(\alu/N102 ), .I1(\alu/N211 ), .S(n5947), .Z(
        \U3/U26/Z_10 ) );
  MUX2D0BWP U4266 ( .I0(\alu/N93 ), .I1(\alu/N202 ), .S(n5947), .Z(
        \U3/U26/Z_1 ) );
  MUX2D0BWP U4267 ( .I0(\alu/N94 ), .I1(\alu/N203 ), .S(n5947), .Z(
        \U3/U26/Z_2 ) );
  MUX2D0BWP U4268 ( .I0(\alu/N95 ), .I1(\alu/N204 ), .S(n5947), .Z(
        \U3/U26/Z_3 ) );
  MUX2D0BWP U4269 ( .I0(\alu/N103 ), .I1(\alu/N212 ), .S(n5947), .Z(
        \U3/U26/Z_11 ) );
  MUX2D0BWP U4270 ( .I0(\alu/N104 ), .I1(\alu/N213 ), .S(n5947), .Z(
        \U3/U26/Z_12 ) );
  MUX2D0BWP U4271 ( .I0(\alu/N105 ), .I1(\alu/N214 ), .S(n5947), .Z(
        \U3/U26/Z_13 ) );
  MUX2D0BWP U4272 ( .I0(\alu/N96 ), .I1(\alu/N205 ), .S(n5947), .Z(
        \U3/U26/Z_4 ) );
  MUX2D0BWP U4273 ( .I0(\alu/N100 ), .I1(\alu/N209 ), .S(n5947), .Z(
        \U3/U26/Z_8 ) );
  MUX2D0BWP U4274 ( .I0(\alu/N99 ), .I1(\alu/N208 ), .S(n5947), .Z(
        \U3/U26/Z_7 ) );
  MUX2D0BWP U4275 ( .I0(\alu/N98 ), .I1(\alu/N207 ), .S(n5947), .Z(
        \U3/U26/Z_6 ) );
  MUX2D0BWP U4276 ( .I0(\alu/N97 ), .I1(\alu/N206 ), .S(n5947), .Z(
        \U3/U26/Z_5 ) );
  MUX2D0BWP U4277 ( .I0(N1182), .I1(N1291), .S(n5987), .Z(\U3/U7/Z_9 ) );
  MUX2D0BWP U4278 ( .I0(N1183), .I1(N1292), .S(n5987), .Z(\U3/U7/Z_10 ) );
  MUX2D0BWP U4279 ( .I0(N1175), .I1(N1284), .S(n5987), .Z(\U3/U7/Z_2 ) );
  MUX2D0BWP U4280 ( .I0(N1176), .I1(N1285), .S(n5987), .Z(\U3/U7/Z_3 ) );
  MUX2D0BWP U4281 ( .I0(N1174), .I1(N1283), .S(n5987), .Z(\U3/U7/Z_1 ) );
  MUX2D0BWP U4282 ( .I0(N1184), .I1(N1293), .S(n5987), .Z(\U3/U7/Z_11 ) );
  MUX2D0BWP U4283 ( .I0(N1177), .I1(N1286), .S(n5987), .Z(\U3/U7/Z_4 ) );
  MUX2D0BWP U4284 ( .I0(N1181), .I1(N1290), .S(n5987), .Z(\U3/U7/Z_8 ) );
  MUX2D0BWP U4285 ( .I0(N1180), .I1(N1289), .S(n5987), .Z(\U3/U7/Z_7 ) );
  MUX2D0BWP U4286 ( .I0(N1185), .I1(N1294), .S(n5987), .Z(\U3/U7/Z_12 ) );
  MUX2D0BWP U4287 ( .I0(N1179), .I1(N1288), .S(n5987), .Z(\U3/U7/Z_6 ) );
  MUX2D0BWP U4288 ( .I0(N1178), .I1(N1287), .S(n5987), .Z(\U3/U7/Z_5 ) );
  MUX2D0BWP U4289 ( .I0(N1186), .I1(N1295), .S(n5987), .Z(\U3/U7/Z_13 ) );
  MUX2D0BWP U4290 ( .I0(\alu/N117 ), .I1(\alu/N226 ), .S(n5947), .Z(
        \U3/U26/Z_25 ) );
  MUX2D0BWP U4291 ( .I0(\alu/N114 ), .I1(\alu/N223 ), .S(n5947), .Z(
        \U3/U26/Z_22 ) );
  MUX2D0BWP U4292 ( .I0(\alu/N113 ), .I1(\alu/N222 ), .S(n5947), .Z(
        \U3/U26/Z_21 ) );
  MUX2D0BWP U4293 ( .I0(\alu/N109 ), .I1(\alu/N218 ), .S(n5947), .Z(
        \U3/U26/Z_17 ) );
  MUX2D0BWP U4294 ( .I0(\alu/N115 ), .I1(\alu/N224 ), .S(n5947), .Z(
        \U3/U26/Z_23 ) );
  MUX2D0BWP U4295 ( .I0(\alu/N116 ), .I1(\alu/N225 ), .S(n5947), .Z(
        \U3/U26/Z_24 ) );
  MUX2D0BWP U4296 ( .I0(\alu/N112 ), .I1(\alu/N221 ), .S(n5947), .Z(
        \U3/U26/Z_20 ) );
  MUX2D0BWP U4297 ( .I0(\alu/N111 ), .I1(\alu/N220 ), .S(n5947), .Z(
        \U3/U26/Z_19 ) );
  MUX2D0BWP U4298 ( .I0(\alu/N110 ), .I1(\alu/N219 ), .S(n5947), .Z(
        \U3/U26/Z_18 ) );
  MUX2D0BWP U4299 ( .I0(N1197), .I1(N1306), .S(n5987), .Z(\U3/U7/Z_24 ) );
  MUX2D0BWP U4300 ( .I0(N1196), .I1(N1305), .S(n5987), .Z(\U3/U7/Z_23 ) );
  MUX2D0BWP U4301 ( .I0(N1195), .I1(N1304), .S(n5987), .Z(\U3/U7/Z_22 ) );
  MUX2D0BWP U4302 ( .I0(N1189), .I1(N1298), .S(n5987), .Z(\U3/U7/Z_16 ) );
  MUX2D0BWP U4303 ( .I0(N1194), .I1(N1303), .S(n5987), .Z(\U3/U7/Z_21 ) );
  MUX2D0BWP U4304 ( .I0(N1193), .I1(N1302), .S(n5987), .Z(\U3/U7/Z_20 ) );
  MUX2D0BWP U4305 ( .I0(N1190), .I1(N1299), .S(n5987), .Z(\U3/U7/Z_17 ) );
  MUX2D0BWP U4306 ( .I0(N1192), .I1(N1301), .S(n5987), .Z(\U3/U7/Z_19 ) );
  MUX2D0BWP U4307 ( .I0(N1191), .I1(N1300), .S(n5987), .Z(\U3/U7/Z_18 ) );
  MUX2D0BWP U4308 ( .I0(\alu/N92 ), .I1(\alu/N201 ), .S(n5947), .Z(
        \U3/U26/Z_0 ) );
  MUX2D0BWP U4309 ( .I0(N1173), .I1(N1282), .S(n5987), .Z(\U3/U7/Z_0 ) );
  MUX2D0BWP U4310 ( .I0(N1198), .I1(N1307), .S(n5987), .Z(\U3/U7/Z_25 ) );
  OR2XD1BWP U4311 ( .A1(n3266), .A2(Reset), .Z(n6180) );
  ND4D1BWP U4312 ( .A1(state[2]), .A2(n7038), .A3(n7436), .A4(n5544), .ZN(
        n7022) );
  INVD1BWP U4313 ( .I(\srf/N15 ), .ZN(n7437) );
  ND4D1BWP U4314 ( .A1(n5867), .A2(cycles[3]), .A3(n5869), .A4(n5873), .ZN(
        n5596) );
  NR2XD0BWP U4315 ( .A1(n7011), .A2(cycles[4]), .ZN(n5600) );
  MUX2D0BWP U4316 ( .I0(\alu/N108 ), .I1(\alu/N217 ), .S(n5947), .Z(
        \U3/U26/Z_16 ) );
  MUX3ND0BWP U4317 ( .I0(n5431), .I1(n5432), .I2(n5433), .S0(func[2]), .S1(
        func[1]), .ZN(result[6]) );
  MUX3ND0BWP U4318 ( .I0(n5435), .I1(n5436), .I2(n5437), .S0(func[2]), .S1(
        func[1]), .ZN(result[7]) );
  MUX3ND0BWP U4319 ( .I0(n5439), .I1(n5440), .I2(n5441), .S0(func[2]), .S1(
        func[1]), .ZN(result[8]) );
  MUX3ND0BWP U4320 ( .I0(n5443), .I1(n5444), .I2(n5445), .S0(func[2]), .S1(
        func[1]), .ZN(result[9]) );
  MUX3ND0BWP U4321 ( .I0(n5427), .I1(n5428), .I2(n5429), .S0(func[2]), .S1(
        func[1]), .ZN(result[5]) );
  MUX3ND0BWP U4322 ( .I0(n5423), .I1(n5424), .I2(n5425), .S0(func[2]), .S1(
        func[1]), .ZN(result[4]) );
  MUX3ND0BWP U4323 ( .I0(n5419), .I1(n5420), .I2(n5421), .S0(func[2]), .S1(
        func[1]), .ZN(result[3]) );
  MUX3ND0BWP U4324 ( .I0(n5407), .I1(n5408), .I2(n5409), .S0(func[2]), .S1(
        func[1]), .ZN(result[0]) );
  MUX3ND0BWP U4325 ( .I0(n5415), .I1(n5416), .I2(n5417), .S0(func[2]), .S1(
        func[1]), .ZN(result[2]) );
  MUX3ND0BWP U4326 ( .I0(n5411), .I1(n5412), .I2(n5413), .S0(func[2]), .S1(
        func[1]), .ZN(result[1]) );
  CKBD1BWP U4327 ( .I(n4681), .Z(n4678) );
  CKBD1BWP U4328 ( .I(n4744), .Z(n4739) );
  CKBD1BWP U4329 ( .I(n4744), .Z(n4738) );
  CKBD1BWP U4330 ( .I(n4744), .Z(n4737) );
  CKBD1BWP U4331 ( .I(n4745), .Z(n4736) );
  CKBD1BWP U4332 ( .I(n4745), .Z(n4735) );
  CKBD1BWP U4333 ( .I(n4745), .Z(n4734) );
  CKBD1BWP U4334 ( .I(n4746), .Z(n4733) );
  CKBD1BWP U4335 ( .I(n4746), .Z(n4732) );
  CKBD1BWP U4336 ( .I(n4746), .Z(n4731) );
  CKBD1BWP U4337 ( .I(n4747), .Z(n4730) );
  CKBD1BWP U4338 ( .I(n4747), .Z(n4729) );
  CKBD1BWP U4339 ( .I(n4747), .Z(n4728) );
  CKBD1BWP U4340 ( .I(n4748), .Z(n4727) );
  CKBD1BWP U4341 ( .I(n4748), .Z(n4726) );
  CKBD1BWP U4342 ( .I(n4748), .Z(n4725) );
  CKBD1BWP U4343 ( .I(n4681), .Z(n4679) );
  CKBD1BWP U4344 ( .I(n4687), .Z(n4660) );
  CKBD1BWP U4345 ( .I(n4687), .Z(n4661) );
  CKBD1BWP U4346 ( .I(n4687), .Z(n4662) );
  CKBD1BWP U4347 ( .I(n4686), .Z(n4663) );
  CKBD1BWP U4348 ( .I(n4686), .Z(n4664) );
  CKBD1BWP U4349 ( .I(n4686), .Z(n4665) );
  CKBD1BWP U4350 ( .I(n4685), .Z(n4666) );
  CKBD1BWP U4351 ( .I(n4685), .Z(n4667) );
  CKBD1BWP U4352 ( .I(n4685), .Z(n4668) );
  CKBD1BWP U4353 ( .I(n4684), .Z(n4669) );
  CKBD1BWP U4354 ( .I(n4684), .Z(n4670) );
  CKBD1BWP U4355 ( .I(n4684), .Z(n4671) );
  CKBD1BWP U4356 ( .I(n4683), .Z(n4672) );
  CKBD1BWP U4357 ( .I(n4683), .Z(n4673) );
  CKBD1BWP U4358 ( .I(n4683), .Z(n4674) );
  CKBD1BWP U4359 ( .I(n4682), .Z(n4675) );
  CKBD1BWP U4360 ( .I(n4682), .Z(n4676) );
  CKBD1BWP U4361 ( .I(n4682), .Z(n4677) );
  CKBD1BWP U4362 ( .I(n4749), .Z(n4724) );
  CKBD1BWP U4363 ( .I(n4749), .Z(n4723) );
  CKBD1BWP U4364 ( .I(n4681), .Z(n4680) );
  CKBD1BWP U4365 ( .I(n4983), .Z(n4946) );
  CKBD1BWP U4366 ( .I(n4987), .Z(n4932) );
  CKBD1BWP U4367 ( .I(n4982), .Z(n4948) );
  CKBD1BWP U4368 ( .I(n4978), .Z(n4959) );
  CKBD1BWP U4369 ( .I(n4979), .Z(n4958) );
  CKBD1BWP U4370 ( .I(n4988), .Z(n4931) );
  CKBD1BWP U4371 ( .I(n4982), .Z(n4947) );
  CKBD1BWP U4372 ( .I(n4975), .Z(n4970) );
  CKBD1BWP U4373 ( .I(n4988), .Z(n4929) );
  CKBD1BWP U4374 ( .I(n4988), .Z(n4930) );
  CKBD1BWP U4375 ( .I(n4980), .Z(n4954) );
  CKBD1BWP U4376 ( .I(n4985), .Z(n4940) );
  CKBD1BWP U4377 ( .I(n4977), .Z(n4964) );
  CKBD1BWP U4378 ( .I(n4979), .Z(n4956) );
  CKBD1BWP U4379 ( .I(n4984), .Z(n4943) );
  CKBD1BWP U4380 ( .I(n4977), .Z(n4962) );
  CKBD1BWP U4381 ( .I(n4979), .Z(n4957) );
  CKBD1BWP U4382 ( .I(n4985), .Z(n4938) );
  CKBD1BWP U4383 ( .I(n4986), .Z(n4935) );
  CKBD1BWP U4384 ( .I(n4984), .Z(n4941) );
  CKBD1BWP U4385 ( .I(n4987), .Z(n4933) );
  CKBD1BWP U4386 ( .I(n4983), .Z(n4944) );
  CKBD1BWP U4387 ( .I(n4978), .Z(n4960) );
  CKBD1BWP U4388 ( .I(n4986), .Z(n4936) );
  CKBD1BWP U4389 ( .I(n4984), .Z(n4942) );
  CKBD1BWP U4390 ( .I(n4985), .Z(n4939) );
  CKBD1BWP U4391 ( .I(n4983), .Z(n4945) );
  CKBD1BWP U4392 ( .I(n4977), .Z(n4963) );
  CKBD1BWP U4393 ( .I(n4978), .Z(n4961) );
  CKBD1BWP U4394 ( .I(n4980), .Z(n4955) );
  CKBD1BWP U4395 ( .I(n4986), .Z(n4937) );
  CKBD1BWP U4396 ( .I(n4987), .Z(n4934) );
  CKBD1BWP U4397 ( .I(n4982), .Z(n4949) );
  CKBD1BWP U4398 ( .I(n4976), .Z(n4965) );
  CKBD1BWP U4399 ( .I(n4981), .Z(n4952) );
  CKBD1BWP U4400 ( .I(n4975), .Z(n4968) );
  CKBD1BWP U4401 ( .I(n4981), .Z(n4950) );
  CKBD1BWP U4402 ( .I(n4976), .Z(n4966) );
  CKBD1BWP U4403 ( .I(n4980), .Z(n4953) );
  CKBD1BWP U4404 ( .I(n4975), .Z(n4969) );
  CKBD1BWP U4405 ( .I(n4981), .Z(n4951) );
  CKBD1BWP U4406 ( .I(n4976), .Z(n4967) );
  CKBD1BWP U4407 ( .I(n5053), .Z(n5016) );
  CKBD1BWP U4408 ( .I(n5057), .Z(n5002) );
  CKBD1BWP U4409 ( .I(n5052), .Z(n5018) );
  CKBD1BWP U4410 ( .I(n5048), .Z(n5029) );
  CKBD1BWP U4411 ( .I(n5049), .Z(n5028) );
  CKBD1BWP U4412 ( .I(n5058), .Z(n5001) );
  CKBD1BWP U4413 ( .I(n5052), .Z(n5017) );
  CKBD1BWP U4414 ( .I(n5045), .Z(n5040) );
  CKBD1BWP U4415 ( .I(n5058), .Z(n4999) );
  CKBD1BWP U4416 ( .I(n5058), .Z(n5000) );
  CKBD1BWP U4417 ( .I(n5050), .Z(n5024) );
  CKBD1BWP U4418 ( .I(n5055), .Z(n5010) );
  CKBD1BWP U4419 ( .I(n5047), .Z(n5034) );
  CKBD1BWP U4420 ( .I(n5049), .Z(n5026) );
  CKBD1BWP U4421 ( .I(n5054), .Z(n5013) );
  CKBD1BWP U4422 ( .I(n5047), .Z(n5032) );
  CKBD1BWP U4423 ( .I(n5049), .Z(n5027) );
  CKBD1BWP U4424 ( .I(n5055), .Z(n5008) );
  CKBD1BWP U4425 ( .I(n5056), .Z(n5005) );
  CKBD1BWP U4426 ( .I(n5054), .Z(n5011) );
  CKBD1BWP U4427 ( .I(n5057), .Z(n5003) );
  CKBD1BWP U4428 ( .I(n5053), .Z(n5014) );
  CKBD1BWP U4429 ( .I(n5048), .Z(n5030) );
  CKBD1BWP U4430 ( .I(n5056), .Z(n5006) );
  CKBD1BWP U4431 ( .I(n5054), .Z(n5012) );
  CKBD1BWP U4432 ( .I(n5055), .Z(n5009) );
  CKBD1BWP U4433 ( .I(n5053), .Z(n5015) );
  CKBD1BWP U4434 ( .I(n5047), .Z(n5033) );
  CKBD1BWP U4435 ( .I(n5048), .Z(n5031) );
  CKBD1BWP U4436 ( .I(n5050), .Z(n5025) );
  CKBD1BWP U4437 ( .I(n5056), .Z(n5007) );
  CKBD1BWP U4438 ( .I(n5057), .Z(n5004) );
  CKBD1BWP U4439 ( .I(n5052), .Z(n5019) );
  CKBD1BWP U4440 ( .I(n5046), .Z(n5035) );
  CKBD1BWP U4441 ( .I(n5051), .Z(n5022) );
  CKBD1BWP U4442 ( .I(n5045), .Z(n5038) );
  CKBD1BWP U4443 ( .I(n5051), .Z(n5020) );
  CKBD1BWP U4444 ( .I(n5046), .Z(n5036) );
  CKBD1BWP U4445 ( .I(n5050), .Z(n5023) );
  CKBD1BWP U4446 ( .I(n5045), .Z(n5039) );
  CKBD1BWP U4447 ( .I(n5051), .Z(n5021) );
  CKBD1BWP U4448 ( .I(n5046), .Z(n5037) );
  CKBD1BWP U4449 ( .I(n4751), .Z(n4744) );
  CKBD1BWP U4450 ( .I(n4751), .Z(n4745) );
  CKBD1BWP U4451 ( .I(n4751), .Z(n4746) );
  CKBD1BWP U4452 ( .I(n4750), .Z(n4747) );
  CKBD1BWP U4453 ( .I(n4750), .Z(n4748) );
  CKBD1BWP U4454 ( .I(n4689), .Z(n4687) );
  CKBD1BWP U4455 ( .I(n4689), .Z(n4686) );
  CKBD1BWP U4456 ( .I(n4690), .Z(n4685) );
  CKBD1BWP U4457 ( .I(n4690), .Z(n4684) );
  CKBD1BWP U4458 ( .I(n4690), .Z(n4683) );
  CKBD1BWP U4459 ( .I(n4691), .Z(n4681) );
  CKBD1BWP U4460 ( .I(n4691), .Z(n4682) );
  CKBD1BWP U4461 ( .I(n4750), .Z(n4749) );
  CKBD1BWP U4462 ( .I(n4743), .Z(n4741) );
  CKBD1BWP U4463 ( .I(n4743), .Z(n4740) );
  CKBD1BWP U4464 ( .I(n4688), .Z(n4659) );
  CKBD1BWP U4465 ( .I(n4689), .Z(n4688) );
  CKBD1BWP U4466 ( .I(n4743), .Z(n4742) );
  CKBD1BWP U4467 ( .I(n4809), .Z(n4768) );
  CKBD1BWP U4468 ( .I(n4811), .Z(n4760) );
  CKBD1BWP U4469 ( .I(n4812), .Z(n4757) );
  CKBD1BWP U4470 ( .I(n4804), .Z(n4781) );
  CKBD1BWP U4471 ( .I(n4813), .Z(n4755) );
  CKBD1BWP U4472 ( .I(n4805), .Z(n4779) );
  CKBD1BWP U4473 ( .I(n4808), .Z(n4770) );
  CKBD1BWP U4474 ( .I(n4805), .Z(n4778) );
  CKBD1BWP U4475 ( .I(n4809), .Z(n4766) );
  CKBD1BWP U4476 ( .I(n4812), .Z(n4758) );
  CKBD1BWP U4477 ( .I(n4809), .Z(n4767) );
  CKBD1BWP U4478 ( .I(n4808), .Z(n4769) );
  CKBD1BWP U4479 ( .I(n4813), .Z(n4756) );
  CKBD1BWP U4480 ( .I(n4812), .Z(n4759) );
  CKBD1BWP U4481 ( .I(n4806), .Z(n4777) );
  CKBD1BWP U4482 ( .I(n4805), .Z(n4780) );
  CKBD1BWP U4483 ( .I(n4801), .Z(n4792) );
  CKBD1BWP U4484 ( .I(n4806), .Z(n4776) );
  CKBD1BWP U4485 ( .I(n4803), .Z(n4784) );
  CKBD1BWP U4486 ( .I(n4802), .Z(n4789) );
  CKBD1BWP U4487 ( .I(n4807), .Z(n4773) );
  CKBD1BWP U4488 ( .I(n4810), .Z(n4765) );
  CKBD1BWP U4489 ( .I(n4802), .Z(n4787) );
  CKBD1BWP U4490 ( .I(n4808), .Z(n4771) );
  CKBD1BWP U4491 ( .I(n4810), .Z(n4763) );
  CKBD1BWP U4492 ( .I(n4800), .Z(n4794) );
  CKBD1BWP U4493 ( .I(n4811), .Z(n4762) );
  CKBD1BWP U4494 ( .I(n4803), .Z(n4786) );
  CKBD1BWP U4495 ( .I(n4801), .Z(n4790) );
  CKBD1BWP U4496 ( .I(n4807), .Z(n4774) );
  CKBD1BWP U4497 ( .I(n4804), .Z(n4782) );
  CKBD1BWP U4498 ( .I(n4801), .Z(n4791) );
  CKBD1BWP U4499 ( .I(n4802), .Z(n4788) );
  CKBD1BWP U4500 ( .I(n4800), .Z(n4793) );
  CKBD1BWP U4501 ( .I(n4806), .Z(n4775) );
  CKBD1BWP U4502 ( .I(n4807), .Z(n4772) );
  CKBD1BWP U4503 ( .I(n4810), .Z(n4764) );
  CKBD1BWP U4504 ( .I(n4811), .Z(n4761) );
  CKBD1BWP U4505 ( .I(n4803), .Z(n4785) );
  CKBD1BWP U4506 ( .I(n4804), .Z(n4783) );
  CKBD1BWP U4507 ( .I(n4800), .Z(n4795) );
  CKBD1BWP U4508 ( .I(n4813), .Z(n4754) );
  CKBD1BWP U4509 ( .I(n4974), .Z(n4971) );
  CKBD1BWP U4510 ( .I(n4974), .Z(n4972) );
  CKBD1BWP U4511 ( .I(n6203), .Z(n4751) );
  CKBD1BWP U4512 ( .I(n6203), .Z(n4750) );
  CKBD1BWP U4513 ( .I(n4989), .Z(n4928) );
  CKBD1BWP U4514 ( .I(n4990), .Z(n4989) );
  CKBD1BWP U4515 ( .I(n4879), .Z(n4838) );
  CKBD1BWP U4516 ( .I(n4881), .Z(n4830) );
  CKBD1BWP U4517 ( .I(n4882), .Z(n4827) );
  CKBD1BWP U4518 ( .I(n4874), .Z(n4851) );
  CKBD1BWP U4519 ( .I(n4883), .Z(n4825) );
  CKBD1BWP U4520 ( .I(n4875), .Z(n4849) );
  CKBD1BWP U4521 ( .I(n4878), .Z(n4840) );
  CKBD1BWP U4522 ( .I(n4875), .Z(n4848) );
  CKBD1BWP U4523 ( .I(n4879), .Z(n4836) );
  CKBD1BWP U4524 ( .I(n4882), .Z(n4828) );
  CKBD1BWP U4525 ( .I(n4879), .Z(n4837) );
  CKBD1BWP U4526 ( .I(n4878), .Z(n4839) );
  CKBD1BWP U4527 ( .I(n4883), .Z(n4826) );
  CKBD1BWP U4528 ( .I(n4882), .Z(n4829) );
  CKBD1BWP U4529 ( .I(n4876), .Z(n4847) );
  CKBD1BWP U4530 ( .I(n4875), .Z(n4850) );
  CKBD1BWP U4531 ( .I(n4871), .Z(n4862) );
  CKBD1BWP U4532 ( .I(n4876), .Z(n4846) );
  CKBD1BWP U4533 ( .I(n4873), .Z(n4854) );
  CKBD1BWP U4534 ( .I(n4872), .Z(n4859) );
  CKBD1BWP U4535 ( .I(n4877), .Z(n4843) );
  CKBD1BWP U4536 ( .I(n4880), .Z(n4835) );
  CKBD1BWP U4537 ( .I(n4872), .Z(n4857) );
  CKBD1BWP U4538 ( .I(n4878), .Z(n4841) );
  CKBD1BWP U4539 ( .I(n4880), .Z(n4833) );
  CKBD1BWP U4540 ( .I(n4870), .Z(n4864) );
  CKBD1BWP U4541 ( .I(n4881), .Z(n4832) );
  CKBD1BWP U4542 ( .I(n4873), .Z(n4856) );
  CKBD1BWP U4543 ( .I(n4871), .Z(n4860) );
  CKBD1BWP U4544 ( .I(n4877), .Z(n4844) );
  CKBD1BWP U4545 ( .I(n4874), .Z(n4852) );
  CKBD1BWP U4546 ( .I(n4871), .Z(n4861) );
  CKBD1BWP U4547 ( .I(n4872), .Z(n4858) );
  CKBD1BWP U4548 ( .I(n4870), .Z(n4863) );
  CKBD1BWP U4549 ( .I(n4876), .Z(n4845) );
  CKBD1BWP U4550 ( .I(n4877), .Z(n4842) );
  CKBD1BWP U4551 ( .I(n4880), .Z(n4834) );
  CKBD1BWP U4552 ( .I(n4881), .Z(n4831) );
  CKBD1BWP U4553 ( .I(n4873), .Z(n4855) );
  CKBD1BWP U4554 ( .I(n4874), .Z(n4853) );
  CKBD1BWP U4555 ( .I(n4870), .Z(n4865) );
  CKBD1BWP U4556 ( .I(n4883), .Z(n4824) );
  CKBD1BWP U4557 ( .I(n5044), .Z(n5041) );
  CKBD1BWP U4558 ( .I(n5044), .Z(n5042) );
  CKBD1BWP U4559 ( .I(n5059), .Z(n4998) );
  CKBD1BWP U4560 ( .I(n5060), .Z(n5059) );
  CKBD1BWP U4561 ( .I(n5093), .Z(n5083) );
  CKBD1BWP U4562 ( .I(n5095), .Z(n5077) );
  CKBD1BWP U4563 ( .I(n5093), .Z(n5082) );
  CKBD1BWP U4564 ( .I(n5096), .Z(n5074) );
  CKBD1BWP U4565 ( .I(n5097), .Z(n5070) );
  CKBD1BWP U4566 ( .I(n5096), .Z(n5075) );
  CKBD1BWP U4567 ( .I(n5096), .Z(n5073) );
  CKBD1BWP U4568 ( .I(n5095), .Z(n5076) );
  CKBD1BWP U4569 ( .I(n5093), .Z(n5084) );
  CKBD1BWP U4570 ( .I(n5094), .Z(n5081) );
  CKBD1BWP U4571 ( .I(n5097), .Z(n5072) );
  CKBD1BWP U4572 ( .I(n5097), .Z(n5071) );
  CKBD1BWP U4573 ( .I(n5095), .Z(n5078) );
  CKBD1BWP U4574 ( .I(n5094), .Z(n5080) );
  CKBD1BWP U4575 ( .I(n5094), .Z(n5079) );
  CKBD1BWP U4576 ( .I(n5091), .Z(n5089) );
  CKBD1BWP U4577 ( .I(n5092), .Z(n5085) );
  CKBD1BWP U4578 ( .I(n5092), .Z(n5086) );
  CKBD1BWP U4579 ( .I(n5091), .Z(n5088) );
  CKBD1BWP U4580 ( .I(n5092), .Z(n5087) );
  CKBD1BWP U4581 ( .I(n5098), .Z(n5069) );
  CKBD1BWP U4582 ( .I(n5098), .Z(n5068) );
  CKBD1BWP U4583 ( .I(n4752), .Z(n4743) );
  CKBD1BWP U4584 ( .I(n6203), .Z(n4752) );
  CKBD1BWP U4585 ( .I(n4692), .Z(n4689) );
  CKBD1BWP U4586 ( .I(n4692), .Z(n4690) );
  CKBD1BWP U4587 ( .I(n4990), .Z(n4987) );
  CKBD1BWP U4588 ( .I(n5060), .Z(n5057) );
  CKBD1BWP U4589 ( .I(n4993), .Z(n4978) );
  CKBD1BWP U4590 ( .I(n5063), .Z(n5048) );
  CKBD1BWP U4591 ( .I(n4992), .Z(n4982) );
  CKBD1BWP U4592 ( .I(n5062), .Z(n5052) );
  CKBD1BWP U4593 ( .I(n4990), .Z(n4988) );
  CKBD1BWP U4594 ( .I(n5060), .Z(n5058) );
  CKBD1BWP U4595 ( .I(n4993), .Z(n4979) );
  CKBD1BWP U4596 ( .I(n5063), .Z(n5049) );
  CKBD1BWP U4597 ( .I(n4991), .Z(n4984) );
  CKBD1BWP U4598 ( .I(n5061), .Z(n5054) );
  CKBD1BWP U4599 ( .I(n4991), .Z(n4985) );
  CKBD1BWP U4600 ( .I(n5061), .Z(n5055) );
  CKBD1BWP U4601 ( .I(n4992), .Z(n4983) );
  CKBD1BWP U4602 ( .I(n5062), .Z(n5053) );
  CKBD1BWP U4603 ( .I(n4994), .Z(n4977) );
  CKBD1BWP U4604 ( .I(n5064), .Z(n5047) );
  CKBD1BWP U4605 ( .I(n4993), .Z(n4980) );
  CKBD1BWP U4606 ( .I(n5063), .Z(n5050) );
  CKBD1BWP U4607 ( .I(n4991), .Z(n4986) );
  CKBD1BWP U4608 ( .I(n5061), .Z(n5056) );
  CKBD1BWP U4609 ( .I(n4994), .Z(n4975) );
  CKBD1BWP U4610 ( .I(n5064), .Z(n5045) );
  CKBD1BWP U4611 ( .I(n4992), .Z(n4981) );
  CKBD1BWP U4612 ( .I(n5062), .Z(n5051) );
  CKBD1BWP U4613 ( .I(n4994), .Z(n4976) );
  CKBD1BWP U4614 ( .I(n5064), .Z(n5046) );
  CKBD1BWP U4615 ( .I(n5091), .Z(n5090) );
  CKBD1BWP U4616 ( .I(n5365), .Z(n5356) );
  CKBD1BWP U4617 ( .I(n5365), .Z(n5355) );
  CKBD1BWP U4618 ( .I(n5365), .Z(n5354) );
  CKBD1BWP U4619 ( .I(n5366), .Z(n5353) );
  CKBD1BWP U4620 ( .I(n5366), .Z(n5352) );
  CKBD1BWP U4621 ( .I(n5367), .Z(n5349) );
  CKBD1BWP U4622 ( .I(n5367), .Z(n5350) );
  CKBD1BWP U4623 ( .I(n5369), .Z(n5342) );
  CKBD1BWP U4624 ( .I(n5369), .Z(n5343) );
  CKBD1BWP U4625 ( .I(n5369), .Z(n5344) );
  CKBD1BWP U4626 ( .I(n5368), .Z(n5345) );
  CKBD1BWP U4627 ( .I(n5368), .Z(n5346) );
  CKBD1BWP U4628 ( .I(n5368), .Z(n5347) );
  CKBD1BWP U4629 ( .I(n5367), .Z(n5348) );
  CKBD1BWP U4630 ( .I(n5366), .Z(n5351) );
  CKBD1BWP U4631 ( .I(n5331), .Z(n5322) );
  CKBD1BWP U4632 ( .I(n5331), .Z(n5321) );
  CKBD1BWP U4633 ( .I(n5331), .Z(n5320) );
  CKBD1BWP U4634 ( .I(n5332), .Z(n5319) );
  CKBD1BWP U4635 ( .I(n5332), .Z(n5318) );
  CKBD1BWP U4636 ( .I(n5333), .Z(n5315) );
  CKBD1BWP U4637 ( .I(n5333), .Z(n5316) );
  CKBD1BWP U4638 ( .I(n5335), .Z(n5308) );
  CKBD1BWP U4639 ( .I(n5335), .Z(n5309) );
  CKBD1BWP U4640 ( .I(n5335), .Z(n5310) );
  CKBD1BWP U4641 ( .I(n5334), .Z(n5311) );
  CKBD1BWP U4642 ( .I(n5334), .Z(n5312) );
  CKBD1BWP U4643 ( .I(n5334), .Z(n5313) );
  CKBD1BWP U4644 ( .I(n5333), .Z(n5314) );
  CKBD1BWP U4645 ( .I(n5332), .Z(n5317) );
  CKBD1BWP U4646 ( .I(n5297), .Z(n5288) );
  CKBD1BWP U4647 ( .I(n5297), .Z(n5287) );
  CKBD1BWP U4648 ( .I(n5297), .Z(n5286) );
  CKBD1BWP U4649 ( .I(n5298), .Z(n5285) );
  CKBD1BWP U4650 ( .I(n5298), .Z(n5284) );
  CKBD1BWP U4651 ( .I(n5299), .Z(n5281) );
  CKBD1BWP U4652 ( .I(n5299), .Z(n5282) );
  CKBD1BWP U4653 ( .I(n5301), .Z(n5274) );
  CKBD1BWP U4654 ( .I(n5301), .Z(n5275) );
  CKBD1BWP U4655 ( .I(n5301), .Z(n5276) );
  CKBD1BWP U4656 ( .I(n5300), .Z(n5277) );
  CKBD1BWP U4657 ( .I(n5300), .Z(n5278) );
  CKBD1BWP U4658 ( .I(n5300), .Z(n5279) );
  CKBD1BWP U4659 ( .I(n5299), .Z(n5280) );
  CKBD1BWP U4660 ( .I(n5298), .Z(n5283) );
  CKBD1BWP U4661 ( .I(n5263), .Z(n5254) );
  CKBD1BWP U4662 ( .I(n5263), .Z(n5253) );
  CKBD1BWP U4663 ( .I(n5263), .Z(n5252) );
  CKBD1BWP U4664 ( .I(n5264), .Z(n5251) );
  CKBD1BWP U4665 ( .I(n5264), .Z(n5250) );
  CKBD1BWP U4666 ( .I(n5265), .Z(n5247) );
  CKBD1BWP U4667 ( .I(n5265), .Z(n5248) );
  CKBD1BWP U4668 ( .I(n5267), .Z(n5240) );
  CKBD1BWP U4669 ( .I(n5267), .Z(n5241) );
  CKBD1BWP U4670 ( .I(n5267), .Z(n5242) );
  CKBD1BWP U4671 ( .I(n5266), .Z(n5243) );
  CKBD1BWP U4672 ( .I(n5266), .Z(n5244) );
  CKBD1BWP U4673 ( .I(n5266), .Z(n5245) );
  CKBD1BWP U4674 ( .I(n5265), .Z(n5246) );
  CKBD1BWP U4675 ( .I(n5264), .Z(n5249) );
  CKBD1BWP U4676 ( .I(n5229), .Z(n5220) );
  CKBD1BWP U4677 ( .I(n5229), .Z(n5219) );
  CKBD1BWP U4678 ( .I(n5229), .Z(n5218) );
  CKBD1BWP U4679 ( .I(n5230), .Z(n5217) );
  CKBD1BWP U4680 ( .I(n5230), .Z(n5216) );
  CKBD1BWP U4681 ( .I(n5231), .Z(n5213) );
  CKBD1BWP U4682 ( .I(n5231), .Z(n5214) );
  CKBD1BWP U4683 ( .I(n5233), .Z(n5206) );
  CKBD1BWP U4684 ( .I(n5233), .Z(n5207) );
  CKBD1BWP U4685 ( .I(n5233), .Z(n5208) );
  CKBD1BWP U4686 ( .I(n5232), .Z(n5209) );
  CKBD1BWP U4687 ( .I(n5232), .Z(n5210) );
  CKBD1BWP U4688 ( .I(n5232), .Z(n5211) );
  CKBD1BWP U4689 ( .I(n5231), .Z(n5212) );
  CKBD1BWP U4690 ( .I(n5230), .Z(n5215) );
  CKBD1BWP U4691 ( .I(n5161), .Z(n5152) );
  CKBD1BWP U4692 ( .I(n5161), .Z(n5151) );
  CKBD1BWP U4693 ( .I(n5161), .Z(n5150) );
  CKBD1BWP U4694 ( .I(n5162), .Z(n5149) );
  CKBD1BWP U4695 ( .I(n5162), .Z(n5148) );
  CKBD1BWP U4696 ( .I(n5163), .Z(n5145) );
  CKBD1BWP U4697 ( .I(n5163), .Z(n5146) );
  CKBD1BWP U4698 ( .I(n5165), .Z(n5138) );
  CKBD1BWP U4699 ( .I(n5165), .Z(n5139) );
  CKBD1BWP U4700 ( .I(n5165), .Z(n5140) );
  CKBD1BWP U4701 ( .I(n5164), .Z(n5141) );
  CKBD1BWP U4702 ( .I(n5164), .Z(n5142) );
  CKBD1BWP U4703 ( .I(n5164), .Z(n5143) );
  CKBD1BWP U4704 ( .I(n5163), .Z(n5144) );
  CKBD1BWP U4705 ( .I(n5162), .Z(n5147) );
  CKBD1BWP U4706 ( .I(n5195), .Z(n5186) );
  CKBD1BWP U4707 ( .I(n5195), .Z(n5185) );
  CKBD1BWP U4708 ( .I(n5195), .Z(n5184) );
  CKBD1BWP U4709 ( .I(n5196), .Z(n5183) );
  CKBD1BWP U4710 ( .I(n5196), .Z(n5182) );
  CKBD1BWP U4711 ( .I(n5197), .Z(n5179) );
  CKBD1BWP U4712 ( .I(n5197), .Z(n5180) );
  CKBD1BWP U4713 ( .I(n5199), .Z(n5172) );
  CKBD1BWP U4714 ( .I(n5199), .Z(n5173) );
  CKBD1BWP U4715 ( .I(n5199), .Z(n5174) );
  CKBD1BWP U4716 ( .I(n5198), .Z(n5175) );
  CKBD1BWP U4717 ( .I(n5198), .Z(n5176) );
  CKBD1BWP U4718 ( .I(n5198), .Z(n5177) );
  CKBD1BWP U4719 ( .I(n5197), .Z(n5178) );
  CKBD1BWP U4720 ( .I(n5196), .Z(n5181) );
  CKBD1BWP U4721 ( .I(n5127), .Z(n5118) );
  CKBD1BWP U4722 ( .I(n5127), .Z(n5117) );
  CKBD1BWP U4723 ( .I(n5127), .Z(n5116) );
  CKBD1BWP U4724 ( .I(n5128), .Z(n5115) );
  CKBD1BWP U4725 ( .I(n5128), .Z(n5114) );
  CKBD1BWP U4726 ( .I(n5129), .Z(n5111) );
  CKBD1BWP U4727 ( .I(n5129), .Z(n5112) );
  CKBD1BWP U4728 ( .I(n5131), .Z(n5104) );
  CKBD1BWP U4729 ( .I(n5131), .Z(n5105) );
  CKBD1BWP U4730 ( .I(n5131), .Z(n5106) );
  CKBD1BWP U4731 ( .I(n5130), .Z(n5107) );
  CKBD1BWP U4732 ( .I(n5130), .Z(n5108) );
  CKBD1BWP U4733 ( .I(n5130), .Z(n5109) );
  CKBD1BWP U4734 ( .I(n5129), .Z(n5110) );
  CKBD1BWP U4735 ( .I(n5128), .Z(n5113) );
  CKBD1BWP U4736 ( .I(n5363), .Z(n5361) );
  CKBD1BWP U4737 ( .I(n5363), .Z(n5360) );
  CKBD1BWP U4738 ( .I(n5364), .Z(n5359) );
  CKBD1BWP U4739 ( .I(n5364), .Z(n5358) );
  CKBD1BWP U4740 ( .I(n5364), .Z(n5357) );
  CKBD1BWP U4741 ( .I(n5329), .Z(n5327) );
  CKBD1BWP U4742 ( .I(n5329), .Z(n5326) );
  CKBD1BWP U4743 ( .I(n5330), .Z(n5325) );
  CKBD1BWP U4744 ( .I(n5330), .Z(n5324) );
  CKBD1BWP U4745 ( .I(n5330), .Z(n5323) );
  CKBD1BWP U4746 ( .I(n5295), .Z(n5293) );
  CKBD1BWP U4747 ( .I(n5295), .Z(n5292) );
  CKBD1BWP U4748 ( .I(n5296), .Z(n5291) );
  CKBD1BWP U4749 ( .I(n5296), .Z(n5290) );
  CKBD1BWP U4750 ( .I(n5296), .Z(n5289) );
  CKBD1BWP U4751 ( .I(n5261), .Z(n5259) );
  CKBD1BWP U4752 ( .I(n5261), .Z(n5258) );
  CKBD1BWP U4753 ( .I(n5262), .Z(n5257) );
  CKBD1BWP U4754 ( .I(n5262), .Z(n5256) );
  CKBD1BWP U4755 ( .I(n5262), .Z(n5255) );
  CKBD1BWP U4756 ( .I(n5227), .Z(n5225) );
  CKBD1BWP U4757 ( .I(n5227), .Z(n5224) );
  CKBD1BWP U4758 ( .I(n5228), .Z(n5223) );
  CKBD1BWP U4759 ( .I(n5228), .Z(n5222) );
  CKBD1BWP U4760 ( .I(n5228), .Z(n5221) );
  CKBD1BWP U4761 ( .I(n5159), .Z(n5157) );
  CKBD1BWP U4762 ( .I(n5159), .Z(n5156) );
  CKBD1BWP U4763 ( .I(n5160), .Z(n5155) );
  CKBD1BWP U4764 ( .I(n5160), .Z(n5154) );
  CKBD1BWP U4765 ( .I(n5160), .Z(n5153) );
  CKBD1BWP U4766 ( .I(n5193), .Z(n5191) );
  CKBD1BWP U4767 ( .I(n5193), .Z(n5190) );
  CKBD1BWP U4768 ( .I(n5194), .Z(n5189) );
  CKBD1BWP U4769 ( .I(n5194), .Z(n5188) );
  CKBD1BWP U4770 ( .I(n5194), .Z(n5187) );
  CKBD1BWP U4771 ( .I(n5125), .Z(n5123) );
  CKBD1BWP U4772 ( .I(n5125), .Z(n5122) );
  CKBD1BWP U4773 ( .I(n5126), .Z(n5121) );
  CKBD1BWP U4774 ( .I(n5126), .Z(n5120) );
  CKBD1BWP U4775 ( .I(n5126), .Z(n5119) );
  CKBD1BWP U4776 ( .I(n4974), .Z(n4973) );
  CKBD1BWP U4777 ( .I(n5396), .Z(n5391) );
  CKBD1BWP U4778 ( .I(n5396), .Z(n5390) );
  CKBD1BWP U4779 ( .I(n5396), .Z(n5389) );
  CKBD1BWP U4780 ( .I(n5397), .Z(n5388) );
  CKBD1BWP U4781 ( .I(n5397), .Z(n5387) );
  CKBD1BWP U4782 ( .I(n5397), .Z(n5386) );
  CKBD1BWP U4783 ( .I(n5398), .Z(n5385) );
  CKBD1BWP U4784 ( .I(n5399), .Z(n5382) );
  CKBD1BWP U4785 ( .I(n5398), .Z(n5383) );
  CKBD1BWP U4786 ( .I(n5398), .Z(n5384) );
  CKBD1BWP U4787 ( .I(n5400), .Z(n5377) );
  CKBD1BWP U4788 ( .I(n5400), .Z(n5378) );
  CKBD1BWP U4789 ( .I(n5400), .Z(n5379) );
  CKBD1BWP U4790 ( .I(n5399), .Z(n5380) );
  CKBD1BWP U4791 ( .I(n5399), .Z(n5381) );
  CKBD1BWP U4792 ( .I(n5401), .Z(n5375) );
  CKBD1BWP U4793 ( .I(n5401), .Z(n5376) );
  CKBD1BWP U4794 ( .I(n4717), .Z(n4694) );
  CKBD1BWP U4795 ( .I(n4717), .Z(n4695) );
  CKBD1BWP U4796 ( .I(n4717), .Z(n4696) );
  CKBD1BWP U4797 ( .I(n4716), .Z(n4697) );
  CKBD1BWP U4798 ( .I(n4716), .Z(n4698) );
  CKBD1BWP U4799 ( .I(n4716), .Z(n4699) );
  CKBD1BWP U4800 ( .I(n4715), .Z(n4700) );
  CKBD1BWP U4801 ( .I(n4715), .Z(n4701) );
  CKBD1BWP U4802 ( .I(n4715), .Z(n4702) );
  CKBD1BWP U4803 ( .I(n4714), .Z(n4703) );
  CKBD1BWP U4804 ( .I(n4714), .Z(n4704) );
  CKBD1BWP U4805 ( .I(n4714), .Z(n4705) );
  CKBD1BWP U4806 ( .I(n4713), .Z(n4706) );
  CKBD1BWP U4807 ( .I(n4713), .Z(n4707) );
  CKBD1BWP U4808 ( .I(n4713), .Z(n4708) );
  CKBD1BWP U4809 ( .I(n4692), .Z(n4691) );
  CKBD1BWP U4810 ( .I(n4655), .Z(n4630) );
  CKBD1BWP U4811 ( .I(n4654), .Z(n4633) );
  CKBD1BWP U4812 ( .I(n4654), .Z(n4632) );
  CKBD1BWP U4813 ( .I(n4650), .Z(n4645) );
  CKBD1BWP U4814 ( .I(n4650), .Z(n4644) );
  CKBD1BWP U4815 ( .I(n4651), .Z(n4642) );
  CKBD1BWP U4816 ( .I(n4651), .Z(n4641) );
  CKBD1BWP U4817 ( .I(n4651), .Z(n4640) );
  CKBD1BWP U4818 ( .I(n4650), .Z(n4643) );
  CKBD1BWP U4819 ( .I(n4654), .Z(n4631) );
  CKBD1BWP U4820 ( .I(n4652), .Z(n4639) );
  CKBD1BWP U4821 ( .I(n4652), .Z(n4638) );
  CKBD1BWP U4822 ( .I(n4652), .Z(n4637) );
  CKBD1BWP U4823 ( .I(n4653), .Z(n4636) );
  CKBD1BWP U4824 ( .I(n4653), .Z(n4635) );
  CKBD1BWP U4825 ( .I(n4653), .Z(n4634) );
  CKBD1BWP U4826 ( .I(n4655), .Z(n4629) );
  CKBD1BWP U4827 ( .I(n5044), .Z(n5043) );
  CKBD1BWP U4828 ( .I(n5363), .Z(n5362) );
  CKBD1BWP U4829 ( .I(n5295), .Z(n5294) );
  CKBD1BWP U4830 ( .I(n5227), .Z(n5226) );
  CKBD1BWP U4831 ( .I(n5159), .Z(n5158) );
  CKBD1BWP U4832 ( .I(n5329), .Z(n5328) );
  CKBD1BWP U4833 ( .I(n5261), .Z(n5260) );
  CKBD1BWP U4834 ( .I(n5193), .Z(n5192) );
  CKBD1BWP U4835 ( .I(n5125), .Z(n5124) );
  CKBD1BWP U4836 ( .I(n4799), .Z(n4797) );
  CKBD1BWP U4837 ( .I(n4799), .Z(n4796) );
  CKBD1BWP U4838 ( .I(n4814), .Z(n4753) );
  CKBD1BWP U4839 ( .I(n4815), .Z(n4814) );
  CKBD1BWP U4840 ( .I(n6201), .Z(n4692) );
  CKBD1BWP U4841 ( .I(n4869), .Z(n4867) );
  CKBD1BWP U4842 ( .I(n4869), .Z(n4866) );
  CKBD1BWP U4843 ( .I(n4884), .Z(n4823) );
  CKBD1BWP U4844 ( .I(n4885), .Z(n4884) );
  CKBD1BWP U4845 ( .I(n4921), .Z(n4899) );
  CKBD1BWP U4846 ( .I(n4922), .Z(n4895) );
  CKBD1BWP U4847 ( .I(n4921), .Z(n4900) );
  CKBD1BWP U4848 ( .I(n4920), .Z(n4901) );
  CKBD1BWP U4849 ( .I(n4922), .Z(n4896) );
  CKBD1BWP U4850 ( .I(n4919), .Z(n4905) );
  CKBD1BWP U4851 ( .I(n4919), .Z(n4906) );
  CKBD1BWP U4852 ( .I(n4920), .Z(n4903) );
  CKBD1BWP U4853 ( .I(n4918), .Z(n4907) );
  CKBD1BWP U4854 ( .I(n4919), .Z(n4904) );
  CKBD1BWP U4855 ( .I(n4920), .Z(n4902) );
  CKBD1BWP U4856 ( .I(n4921), .Z(n4898) );
  CKBD1BWP U4857 ( .I(n4922), .Z(n4897) );
  CKBD1BWP U4858 ( .I(n4918), .Z(n4909) );
  CKBD1BWP U4859 ( .I(n4918), .Z(n4908) );
  CKBD1BWP U4860 ( .I(n4917), .Z(n4911) );
  CKBD1BWP U4861 ( .I(n4917), .Z(n4912) );
  CKBD1BWP U4862 ( .I(n4917), .Z(n4910) );
  CKBD1BWP U4863 ( .I(n4916), .Z(n4913) );
  CKBD1BWP U4864 ( .I(n4916), .Z(n4914) );
  CKBD1BWP U4865 ( .I(n4923), .Z(n4894) );
  CKBD1BWP U4866 ( .I(n4923), .Z(n4893) );
  CKBD1BWP U4867 ( .I(n4997), .Z(n4990) );
  CKBD1BWP U4868 ( .I(n5067), .Z(n5060) );
  CKBD1BWP U4869 ( .I(n4996), .Z(n4993) );
  CKBD1BWP U4870 ( .I(n5066), .Z(n5063) );
  CKBD1BWP U4871 ( .I(n4997), .Z(n4992) );
  CKBD1BWP U4872 ( .I(n5067), .Z(n5062) );
  CKBD1BWP U4873 ( .I(n4997), .Z(n4991) );
  CKBD1BWP U4874 ( .I(n5067), .Z(n5061) );
  CKBD1BWP U4875 ( .I(n4996), .Z(n4994) );
  CKBD1BWP U4876 ( .I(n5066), .Z(n5064) );
  CKBD1BWP U4877 ( .I(n4657), .Z(n4651) );
  CKBD1BWP U4878 ( .I(n4657), .Z(n4650) );
  CKBD1BWP U4879 ( .I(n4656), .Z(n4654) );
  CKBD1BWP U4880 ( .I(n4657), .Z(n4652) );
  CKBD1BWP U4881 ( .I(n4656), .Z(n4653) );
  CKBD1BWP U4882 ( .I(n5372), .Z(n5365) );
  CKBD1BWP U4883 ( .I(n5371), .Z(n5369) );
  CKBD1BWP U4884 ( .I(n5371), .Z(n5368) );
  CKBD1BWP U4885 ( .I(n5372), .Z(n5367) );
  CKBD1BWP U4886 ( .I(n5372), .Z(n5366) );
  CKBD1BWP U4887 ( .I(n5304), .Z(n5297) );
  CKBD1BWP U4888 ( .I(n5303), .Z(n5301) );
  CKBD1BWP U4889 ( .I(n5303), .Z(n5300) );
  CKBD1BWP U4890 ( .I(n5304), .Z(n5299) );
  CKBD1BWP U4891 ( .I(n5304), .Z(n5298) );
  CKBD1BWP U4892 ( .I(n5236), .Z(n5229) );
  CKBD1BWP U4893 ( .I(n5235), .Z(n5233) );
  CKBD1BWP U4894 ( .I(n5235), .Z(n5232) );
  CKBD1BWP U4895 ( .I(n5236), .Z(n5231) );
  CKBD1BWP U4896 ( .I(n5236), .Z(n5230) );
  CKBD1BWP U4897 ( .I(n5168), .Z(n5161) );
  CKBD1BWP U4898 ( .I(n5167), .Z(n5165) );
  CKBD1BWP U4899 ( .I(n5167), .Z(n5164) );
  CKBD1BWP U4900 ( .I(n5168), .Z(n5163) );
  CKBD1BWP U4901 ( .I(n5168), .Z(n5162) );
  CKBD1BWP U4902 ( .I(n5338), .Z(n5331) );
  CKBD1BWP U4903 ( .I(n5337), .Z(n5335) );
  CKBD1BWP U4904 ( .I(n5337), .Z(n5334) );
  CKBD1BWP U4905 ( .I(n5338), .Z(n5333) );
  CKBD1BWP U4906 ( .I(n5338), .Z(n5332) );
  CKBD1BWP U4907 ( .I(n5270), .Z(n5263) );
  CKBD1BWP U4908 ( .I(n5269), .Z(n5267) );
  CKBD1BWP U4909 ( .I(n5269), .Z(n5266) );
  CKBD1BWP U4910 ( .I(n5270), .Z(n5265) );
  CKBD1BWP U4911 ( .I(n5270), .Z(n5264) );
  CKBD1BWP U4912 ( .I(n4816), .Z(n4811) );
  CKBD1BWP U4913 ( .I(n4886), .Z(n4881) );
  CKBD1BWP U4914 ( .I(n4818), .Z(n4804) );
  CKBD1BWP U4915 ( .I(n4888), .Z(n4874) );
  CKBD1BWP U4916 ( .I(n4816), .Z(n4809) );
  CKBD1BWP U4917 ( .I(n4886), .Z(n4879) );
  CKBD1BWP U4918 ( .I(n4817), .Z(n4808) );
  CKBD1BWP U4919 ( .I(n4887), .Z(n4878) );
  CKBD1BWP U4920 ( .I(n4815), .Z(n4813) );
  CKBD1BWP U4921 ( .I(n4885), .Z(n4883) );
  CKBD1BWP U4922 ( .I(n4815), .Z(n4812) );
  CKBD1BWP U4923 ( .I(n4885), .Z(n4882) );
  CKBD1BWP U4924 ( .I(n4818), .Z(n4805) );
  CKBD1BWP U4925 ( .I(n4888), .Z(n4875) );
  CKBD1BWP U4926 ( .I(n4819), .Z(n4801) );
  CKBD1BWP U4927 ( .I(n4889), .Z(n4871) );
  CKBD1BWP U4928 ( .I(n4819), .Z(n4802) );
  CKBD1BWP U4929 ( .I(n4889), .Z(n4872) );
  CKBD1BWP U4930 ( .I(n4819), .Z(n4800) );
  CKBD1BWP U4931 ( .I(n4889), .Z(n4870) );
  CKBD1BWP U4932 ( .I(n4817), .Z(n4806) );
  CKBD1BWP U4933 ( .I(n4887), .Z(n4876) );
  CKBD1BWP U4934 ( .I(n4817), .Z(n4807) );
  CKBD1BWP U4935 ( .I(n4887), .Z(n4877) );
  CKBD1BWP U4936 ( .I(n4816), .Z(n4810) );
  CKBD1BWP U4937 ( .I(n4886), .Z(n4880) );
  CKBD1BWP U4938 ( .I(n4818), .Z(n4803) );
  CKBD1BWP U4939 ( .I(n4888), .Z(n4873) );
  CKBD1BWP U4940 ( .I(n5403), .Z(n5396) );
  CKBD1BWP U4941 ( .I(n5403), .Z(n5397) );
  CKBD1BWP U4942 ( .I(n5403), .Z(n5398) );
  CKBD1BWP U4943 ( .I(n5402), .Z(n5400) );
  CKBD1BWP U4944 ( .I(n5402), .Z(n5399) );
  CKBD1BWP U4945 ( .I(n5202), .Z(n5195) );
  CKBD1BWP U4946 ( .I(n5201), .Z(n5199) );
  CKBD1BWP U4947 ( .I(n5201), .Z(n5198) );
  CKBD1BWP U4948 ( .I(n5202), .Z(n5197) );
  CKBD1BWP U4949 ( .I(n5202), .Z(n5196) );
  CKBD1BWP U4950 ( .I(n5134), .Z(n5127) );
  CKBD1BWP U4951 ( .I(n5133), .Z(n5131) );
  CKBD1BWP U4952 ( .I(n5133), .Z(n5130) );
  CKBD1BWP U4953 ( .I(n5134), .Z(n5129) );
  CKBD1BWP U4954 ( .I(n5134), .Z(n5128) );
  CKBD1BWP U4955 ( .I(n5100), .Z(n5095) );
  CKBD1BWP U4956 ( .I(n5099), .Z(n5096) );
  CKBD1BWP U4957 ( .I(n5100), .Z(n5093) );
  CKBD1BWP U4958 ( .I(n5099), .Z(n5097) );
  CKBD1BWP U4959 ( .I(n5100), .Z(n5094) );
  CKBD1BWP U4960 ( .I(n4719), .Z(n4717) );
  CKBD1BWP U4961 ( .I(n4719), .Z(n4716) );
  CKBD1BWP U4962 ( .I(n4720), .Z(n4715) );
  CKBD1BWP U4963 ( .I(n4720), .Z(n4714) );
  CKBD1BWP U4964 ( .I(n4720), .Z(n4713) );
  CKBD1BWP U4965 ( .I(n5373), .Z(n5364) );
  CKBD1BWP U4966 ( .I(n5373), .Z(n5363) );
  CKBD1BWP U4967 ( .I(n5305), .Z(n5296) );
  CKBD1BWP U4968 ( .I(n5305), .Z(n5295) );
  CKBD1BWP U4969 ( .I(n5237), .Z(n5228) );
  CKBD1BWP U4970 ( .I(n5237), .Z(n5227) );
  CKBD1BWP U4971 ( .I(n5169), .Z(n5160) );
  CKBD1BWP U4972 ( .I(n5169), .Z(n5159) );
  CKBD1BWP U4973 ( .I(n5339), .Z(n5330) );
  CKBD1BWP U4974 ( .I(n5339), .Z(n5329) );
  CKBD1BWP U4975 ( .I(n5271), .Z(n5262) );
  CKBD1BWP U4976 ( .I(n5271), .Z(n5261) );
  CKBD1BWP U4977 ( .I(n5203), .Z(n5194) );
  CKBD1BWP U4978 ( .I(n5203), .Z(n5193) );
  CKBD1BWP U4979 ( .I(n5135), .Z(n5126) );
  CKBD1BWP U4980 ( .I(n5135), .Z(n5125) );
  CKBD1BWP U4981 ( .I(n5101), .Z(n5091) );
  CKBD1BWP U4982 ( .I(n5101), .Z(n5092) );
  CKBD1BWP U4983 ( .I(n4995), .Z(n4974) );
  CKBD1BWP U4984 ( .I(n4996), .Z(n4995) );
  CKBD1BWP U4985 ( .I(n5065), .Z(n5044) );
  CKBD1BWP U4986 ( .I(n5066), .Z(n5065) );
  CKBD1BWP U4987 ( .I(n4916), .Z(n4915) );
  CKBD1BWP U4988 ( .I(n4799), .Z(n4798) );
  CKBD1BWP U4989 ( .I(n5395), .Z(n5393) );
  CKBD1BWP U4990 ( .I(n5395), .Z(n5392) );
  CKBD1BWP U4991 ( .I(n5395), .Z(n5394) );
  CKBD1BWP U4992 ( .I(n5370), .Z(n5341) );
  CKBD1BWP U4993 ( .I(n5371), .Z(n5370) );
  CKBD1BWP U4994 ( .I(n5336), .Z(n5307) );
  CKBD1BWP U4995 ( .I(n5337), .Z(n5336) );
  CKBD1BWP U4996 ( .I(n5302), .Z(n5273) );
  CKBD1BWP U4997 ( .I(n5303), .Z(n5302) );
  CKBD1BWP U4998 ( .I(n5268), .Z(n5239) );
  CKBD1BWP U4999 ( .I(n5269), .Z(n5268) );
  CKBD1BWP U5000 ( .I(n5234), .Z(n5205) );
  CKBD1BWP U5001 ( .I(n5235), .Z(n5234) );
  CKBD1BWP U5002 ( .I(n5166), .Z(n5137) );
  CKBD1BWP U5003 ( .I(n5167), .Z(n5166) );
  CKBD1BWP U5004 ( .I(n5200), .Z(n5171) );
  CKBD1BWP U5005 ( .I(n5201), .Z(n5200) );
  CKBD1BWP U5006 ( .I(n5132), .Z(n5103) );
  CKBD1BWP U5007 ( .I(n5133), .Z(n5132) );
  CKBD1BWP U5008 ( .I(n4712), .Z(n4709) );
  CKBD1BWP U5009 ( .I(n4712), .Z(n4710) );
  CKBD1BWP U5010 ( .I(n4656), .Z(n4655) );
  CKBD1BWP U5011 ( .I(n4718), .Z(n4693) );
  CKBD1BWP U5012 ( .I(n4719), .Z(n4718) );
  CKBD1BWP U5013 ( .I(n5402), .Z(n5401) );
  CKBD1BWP U5014 ( .I(n5099), .Z(n5098) );
  CKBD1BWP U5015 ( .I(n4649), .Z(n4647) );
  CKBD1BWP U5016 ( .I(n4649), .Z(n4646) );
  CKBD1BWP U5017 ( .I(n4649), .Z(n4648) );
  CKBD1BWP U5018 ( .I(n4869), .Z(n4868) );
  CKBD1BWP U5019 ( .I(n4712), .Z(n4711) );
  CKBD1BWP U5020 ( .I(\vrf/N13 ), .Z(n5067) );
  CKBD1BWP U5021 ( .I(\vrf/N13 ), .Z(n5066) );
  CKBD1BWP U5022 ( .I(\vrf/N12 ), .Z(n4997) );
  CKBD1BWP U5023 ( .I(\vrf/N12 ), .Z(n4996) );
  CKBD1BWP U5024 ( .I(n5524), .Z(n4657) );
  CKBD1BWP U5025 ( .I(n5524), .Z(n4656) );
  CKBD1BWP U5026 ( .I(n5374), .Z(n5371) );
  CKBD1BWP U5027 ( .I(n5374), .Z(n5372) );
  CKBD1BWP U5028 ( .I(n5306), .Z(n5303) );
  CKBD1BWP U5029 ( .I(n5306), .Z(n5304) );
  CKBD1BWP U5030 ( .I(n5238), .Z(n5235) );
  CKBD1BWP U5031 ( .I(n5238), .Z(n5236) );
  CKBD1BWP U5032 ( .I(n5170), .Z(n5167) );
  CKBD1BWP U5033 ( .I(n5170), .Z(n5168) );
  CKBD1BWP U5034 ( .I(n5272), .Z(n5269) );
  CKBD1BWP U5035 ( .I(n5272), .Z(n5270) );
  CKBD1BWP U5036 ( .I(n5340), .Z(n5337) );
  CKBD1BWP U5037 ( .I(n5340), .Z(n5338) );
  CKBD1BWP U5038 ( .I(n4822), .Z(n4816) );
  CKBD1BWP U5039 ( .I(n4892), .Z(n4886) );
  CKBD1BWP U5040 ( .I(n4822), .Z(n4815) );
  CKBD1BWP U5041 ( .I(n4892), .Z(n4885) );
  CKBD1BWP U5042 ( .I(n4821), .Z(n4818) );
  CKBD1BWP U5043 ( .I(n4891), .Z(n4888) );
  CKBD1BWP U5044 ( .I(n4821), .Z(n4819) );
  CKBD1BWP U5045 ( .I(n4891), .Z(n4889) );
  CKBD1BWP U5046 ( .I(n4822), .Z(n4817) );
  CKBD1BWP U5047 ( .I(n4892), .Z(n4887) );
  CKBD1BWP U5048 ( .I(n5405), .Z(n5403) );
  CKBD1BWP U5049 ( .I(n5405), .Z(n5402) );
  CKBD1BWP U5050 ( .I(n4658), .Z(n4649) );
  CKBD1BWP U5051 ( .I(n5524), .Z(n4658) );
  CKBD1BWP U5052 ( .I(n5204), .Z(n5201) );
  CKBD1BWP U5053 ( .I(n5204), .Z(n5202) );
  CKBD1BWP U5054 ( .I(n5136), .Z(n5133) );
  CKBD1BWP U5055 ( .I(n5136), .Z(n5134) );
  CKBD1BWP U5056 ( .I(n5102), .Z(n5100) );
  CKBD1BWP U5057 ( .I(n5102), .Z(n5099) );
  CKBD1BWP U5058 ( .I(n4722), .Z(n4719) );
  CKBD1BWP U5059 ( .I(n4722), .Z(n4720) );
  CKBD1BWP U5060 ( .I(n4924), .Z(n4921) );
  CKBD1BWP U5061 ( .I(n4925), .Z(n4920) );
  CKBD1BWP U5062 ( .I(n4924), .Z(n4922) );
  CKBD1BWP U5063 ( .I(n4925), .Z(n4919) );
  CKBD1BWP U5064 ( .I(n4925), .Z(n4918) );
  CKBD1BWP U5065 ( .I(n4926), .Z(n4917) );
  CKBD1BWP U5066 ( .I(n4926), .Z(n4916) );
  CKBD1BWP U5067 ( .I(n4820), .Z(n4799) );
  CKBD1BWP U5068 ( .I(n4821), .Z(n4820) );
  CKBD1BWP U5069 ( .I(n4890), .Z(n4869) );
  CKBD1BWP U5070 ( .I(n4891), .Z(n4890) );
  CKBD1BWP U5071 ( .I(n5404), .Z(n5395) );
  CKBD1BWP U5072 ( .I(n5405), .Z(n5404) );
  CKBD1BWP U5073 ( .I(n4721), .Z(n4712) );
  CKBD1BWP U5074 ( .I(n4722), .Z(n4721) );
  CKBD1BWP U5075 ( .I(n5374), .Z(n5373) );
  CKBD1BWP U5076 ( .I(n5306), .Z(n5305) );
  CKBD1BWP U5077 ( .I(n5238), .Z(n5237) );
  CKBD1BWP U5078 ( .I(n5170), .Z(n5169) );
  CKBD1BWP U5079 ( .I(n5272), .Z(n5271) );
  CKBD1BWP U5080 ( .I(n5340), .Z(n5339) );
  CKBD1BWP U5081 ( .I(n5204), .Z(n5203) );
  CKBD1BWP U5082 ( .I(n5136), .Z(n5135) );
  CKBD1BWP U5083 ( .I(n5102), .Z(n5101) );
  CKBD1BWP U5084 ( .I(n4924), .Z(n4923) );
  CKND0BWP U5085 ( .I(n7437), .ZN(n5498) );
  CKND0BWP U5086 ( .I(n7437), .ZN(n5497) );
  CKND0BWP U5087 ( .I(n7437), .ZN(n5500) );
  CKND0BWP U5088 ( .I(n7437), .ZN(n5499) );
  CKND0BWP U5089 ( .I(n7437), .ZN(n5502) );
  CKND0BWP U5090 ( .I(n7437), .ZN(n5501) );
  CKND0BWP U5091 ( .I(n7437), .ZN(n5504) );
  CKND0BWP U5092 ( .I(n7437), .ZN(n5503) );
  CKND0BWP U5093 ( .I(n7437), .ZN(n5506) );
  CKND0BWP U5094 ( .I(n7437), .ZN(n5505) );
  CKND0BWP U5095 ( .I(n7437), .ZN(n5508) );
  CKND0BWP U5096 ( .I(n7437), .ZN(n5507) );
  CKND0BWP U5097 ( .I(n7437), .ZN(n5510) );
  CKND0BWP U5098 ( .I(n7437), .ZN(n5509) );
  CKND0BWP U5099 ( .I(n7437), .ZN(n5512) );
  CKND0BWP U5100 ( .I(n7437), .ZN(n5511) );
  CKND0BWP U5101 ( .I(n7437), .ZN(n5514) );
  CKND0BWP U5102 ( .I(n7437), .ZN(n5513) );
  CKND0BWP U5103 ( .I(n7437), .ZN(n5516) );
  CKND0BWP U5104 ( .I(n7437), .ZN(n5515) );
  CKND1BWP U5105 ( .I(n7437), .ZN(n5518) );
  CKND1BWP U5106 ( .I(n7437), .ZN(n5517) );
  INVD1BWP U5107 ( .I(n7437), .ZN(n5520) );
  INVD1BWP U5108 ( .I(n7437), .ZN(n5519) );
  INVD1BWP U5109 ( .I(n7437), .ZN(n5522) );
  INVD1BWP U5110 ( .I(n7437), .ZN(n5521) );
  INVD1BWP U5111 ( .I(n7437), .ZN(n5523) );
  INVD1BWP U5112 ( .I(n7438), .ZN(n5486) );
  CKND0BWP U5113 ( .I(n7438), .ZN(n5487) );
  CKND0BWP U5114 ( .I(n7438), .ZN(n5488) );
  CKND0BWP U5115 ( .I(n7438), .ZN(n5489) );
  CKND0BWP U5116 ( .I(n7438), .ZN(n5490) );
  CKND0BWP U5117 ( .I(n7438), .ZN(n5491) );
  CKND0BWP U5118 ( .I(n7438), .ZN(n5492) );
  CKND0BWP U5119 ( .I(n7438), .ZN(n5493) );
  CKND0BWP U5120 ( .I(n7438), .ZN(n5494) );
  CKND0BWP U5121 ( .I(n7438), .ZN(n5495) );
  CKND0BWP U5122 ( .I(n7438), .ZN(n5496) );
  CKBD1BWP U5123 ( .I(\vrf/N296 ), .Z(n5374) );
  CKBD1BWP U5124 ( .I(\vrf/N290 ), .Z(n5306) );
  CKBD1BWP U5125 ( .I(\vrf/N284 ), .Z(n5238) );
  CKBD1BWP U5126 ( .I(\vrf/N278 ), .Z(n5170) );
  CKBD1BWP U5127 ( .I(\vrf/N9 ), .Z(n4822) );
  CKBD1BWP U5128 ( .I(\vrf/N10 ), .Z(n4892) );
  CKBD1BWP U5129 ( .I(\vrf/N9 ), .Z(n4821) );
  CKBD1BWP U5130 ( .I(\vrf/N10 ), .Z(n4891) );
  CKBD1BWP U5131 ( .I(\vrf/N293 ), .Z(n5340) );
  CKBD1BWP U5132 ( .I(\vrf/N287 ), .Z(n5272) );
  CKBD1BWP U5133 ( .I(N4322), .Z(n5405) );
  AN2XD1BWP U5134 ( .A1(\alu/N991 ), .A2(n5485), .Z(n5442) );
  AN2XD1BWP U5135 ( .A1(\alu/N989 ), .A2(n5485), .Z(n5434) );
  AN2XD1BWP U5136 ( .A1(\alu/N988 ), .A2(n5485), .Z(n5430) );
  AN2XD1BWP U5137 ( .A1(\alu/N987 ), .A2(n5485), .Z(n5426) );
  AN2XD1BWP U5138 ( .A1(\alu/N986 ), .A2(n5485), .Z(n5422) );
  AN2XD1BWP U5139 ( .A1(\alu/N985 ), .A2(n5485), .Z(n5418) );
  AN2XD1BWP U5140 ( .A1(\alu/N984 ), .A2(n5485), .Z(n5414) );
  AN2XD1BWP U5141 ( .A1(\alu/N983 ), .A2(n5485), .Z(n5410) );
  AN2XD1BWP U5142 ( .A1(\alu/N990 ), .A2(n5485), .Z(n5438) );
  CKBD1BWP U5143 ( .I(\vrf/N14 ), .Z(n5102) );
  AN2XD1BWP U5144 ( .A1(\alu/N982 ), .A2(n5485), .Z(n5406) );
  CKBD1BWP U5145 ( .I(n6202), .Z(n4722) );
  CKBD1BWP U5146 ( .I(\vrf/N281 ), .Z(n5204) );
  CKBD1BWP U5147 ( .I(\vrf/N217 ), .Z(n5136) );
  AN2XD1BWP U5148 ( .A1(\alu/N835 ), .A2(n5485), .Z(n5458) );
  AN2XD1BWP U5149 ( .A1(\alu/N836 ), .A2(n5485), .Z(n5462) );
  AN2XD1BWP U5150 ( .A1(\alu/N834 ), .A2(n5485), .Z(n5454) );
  AN2XD1BWP U5151 ( .A1(\alu/N999 ), .A2(n5485), .Z(n5446) );
  AN2XD1BWP U5152 ( .A1(\alu/N833 ), .A2(n5485), .Z(n5450) );
  INVD1BWP U5153 ( .I(n5466), .ZN(n5484) );
  CKBD1BWP U5154 ( .I(n4927), .Z(n4924) );
  CKBD1BWP U5155 ( .I(n4927), .Z(n4925) );
  CKBD1BWP U5156 ( .I(n4927), .Z(n4926) );
  MUX2ND0BWP U5157 ( .I0(n3425), .I1(n3426), .S(n5486), .ZN(\srf/N20 ) );
  MUX4ND0BWP U5158 ( .I0(\srf/regTable[0][15] ), .I1(\srf/regTable[1][15] ), 
        .I2(\srf/regTable[2][15] ), .I3(\srf/regTable[3][15] ), .S0(n5497), 
        .S1(\srf/N16 ), .ZN(n3425) );
  MUX4ND0BWP U5159 ( .I0(\srf/regTable[4][15] ), .I1(\srf/regTable[5][15] ), 
        .I2(\srf/regTable[6][15] ), .I3(\srf/regTable[7][15] ), .S0(n5498), 
        .S1(\srf/N16 ), .ZN(n3426) );
  MUX2ND0BWP U5160 ( .I0(n3427), .I1(n3428), .S(n5487), .ZN(\srf/N21 ) );
  MUX4ND0BWP U5161 ( .I0(\srf/regTable[0][14] ), .I1(\srf/regTable[1][14] ), 
        .I2(\srf/regTable[2][14] ), .I3(\srf/regTable[3][14] ), .S0(n5499), 
        .S1(\srf/N16 ), .ZN(n3427) );
  MUX4ND0BWP U5162 ( .I0(\srf/regTable[4][14] ), .I1(\srf/regTable[5][14] ), 
        .I2(\srf/regTable[6][14] ), .I3(\srf/regTable[7][14] ), .S0(n5500), 
        .S1(\srf/N16 ), .ZN(n3428) );
  MUX2ND0BWP U5163 ( .I0(n3429), .I1(n3430), .S(n5488), .ZN(\srf/N22 ) );
  MUX4ND0BWP U5164 ( .I0(\srf/regTable[0][13] ), .I1(\srf/regTable[1][13] ), 
        .I2(\srf/regTable[2][13] ), .I3(\srf/regTable[3][13] ), .S0(n5501), 
        .S1(\srf/N16 ), .ZN(n3429) );
  MUX4ND0BWP U5165 ( .I0(\srf/regTable[4][13] ), .I1(\srf/regTable[5][13] ), 
        .I2(\srf/regTable[6][13] ), .I3(\srf/regTable[7][13] ), .S0(n5502), 
        .S1(\srf/N16 ), .ZN(n3430) );
  MUX2ND0BWP U5166 ( .I0(n3431), .I1(n3432), .S(n5489), .ZN(\srf/N23 ) );
  MUX4ND0BWP U5167 ( .I0(\srf/regTable[0][12] ), .I1(\srf/regTable[1][12] ), 
        .I2(\srf/regTable[2][12] ), .I3(\srf/regTable[3][12] ), .S0(n5503), 
        .S1(\srf/N16 ), .ZN(n3431) );
  MUX4ND0BWP U5168 ( .I0(\srf/regTable[4][12] ), .I1(\srf/regTable[5][12] ), 
        .I2(\srf/regTable[6][12] ), .I3(\srf/regTable[7][12] ), .S0(n5504), 
        .S1(\srf/N16 ), .ZN(n3432) );
  MUX2ND0BWP U5169 ( .I0(n3433), .I1(n3434), .S(n5490), .ZN(\srf/N24 ) );
  MUX4ND0BWP U5170 ( .I0(\srf/regTable[0][11] ), .I1(\srf/regTable[1][11] ), 
        .I2(\srf/regTable[2][11] ), .I3(\srf/regTable[3][11] ), .S0(n5505), 
        .S1(\srf/N16 ), .ZN(n3433) );
  MUX4ND0BWP U5171 ( .I0(\srf/regTable[4][11] ), .I1(\srf/regTable[5][11] ), 
        .I2(\srf/regTable[6][11] ), .I3(\srf/regTable[7][11] ), .S0(n5506), 
        .S1(\srf/N16 ), .ZN(n3434) );
  MUX2ND0BWP U5172 ( .I0(n3435), .I1(n3436), .S(n5491), .ZN(\srf/N25 ) );
  MUX4ND0BWP U5173 ( .I0(\srf/regTable[0][10] ), .I1(\srf/regTable[1][10] ), 
        .I2(\srf/regTable[2][10] ), .I3(\srf/regTable[3][10] ), .S0(n5507), 
        .S1(\srf/N16 ), .ZN(n3435) );
  MUX4ND0BWP U5174 ( .I0(\srf/regTable[4][10] ), .I1(\srf/regTable[5][10] ), 
        .I2(\srf/regTable[6][10] ), .I3(\srf/regTable[7][10] ), .S0(n5508), 
        .S1(\srf/N16 ), .ZN(n3436) );
  MUX2ND0BWP U5175 ( .I0(n3437), .I1(n3438), .S(n5492), .ZN(\srf/N26 ) );
  MUX4ND0BWP U5176 ( .I0(\srf/regTable[0][9] ), .I1(\srf/regTable[1][9] ), 
        .I2(\srf/regTable[2][9] ), .I3(\srf/regTable[3][9] ), .S0(n5509), .S1(
        \srf/N16 ), .ZN(n3437) );
  MUX4ND0BWP U5177 ( .I0(\srf/regTable[4][9] ), .I1(\srf/regTable[5][9] ), 
        .I2(\srf/regTable[6][9] ), .I3(\srf/regTable[7][9] ), .S0(n5510), .S1(
        \srf/N16 ), .ZN(n3438) );
  MUX2ND0BWP U5178 ( .I0(n3439), .I1(n3440), .S(n5493), .ZN(\srf/N27 ) );
  MUX4ND0BWP U5179 ( .I0(\srf/regTable[0][8] ), .I1(\srf/regTable[1][8] ), 
        .I2(\srf/regTable[2][8] ), .I3(\srf/regTable[3][8] ), .S0(n5511), .S1(
        \srf/N16 ), .ZN(n3439) );
  MUX4ND0BWP U5180 ( .I0(\srf/regTable[4][8] ), .I1(\srf/regTable[5][8] ), 
        .I2(\srf/regTable[6][8] ), .I3(\srf/regTable[7][8] ), .S0(n5512), .S1(
        \srf/N16 ), .ZN(n3440) );
  MUX2ND0BWP U5181 ( .I0(n3441), .I1(n3442), .S(n5494), .ZN(\srf/N28 ) );
  MUX4ND0BWP U5182 ( .I0(\srf/regTable[0][7] ), .I1(\srf/regTable[1][7] ), 
        .I2(\srf/regTable[2][7] ), .I3(\srf/regTable[3][7] ), .S0(n5513), .S1(
        \srf/N16 ), .ZN(n3441) );
  MUX4ND0BWP U5183 ( .I0(\srf/regTable[4][7] ), .I1(\srf/regTable[5][7] ), 
        .I2(\srf/regTable[6][7] ), .I3(\srf/regTable[7][7] ), .S0(n5514), .S1(
        \srf/N16 ), .ZN(n3442) );
  MUX2ND0BWP U5184 ( .I0(n3443), .I1(n3444), .S(n5495), .ZN(\srf/N29 ) );
  MUX4ND0BWP U5185 ( .I0(\srf/regTable[0][6] ), .I1(\srf/regTable[1][6] ), 
        .I2(\srf/regTable[2][6] ), .I3(\srf/regTable[3][6] ), .S0(n5515), .S1(
        \srf/N16 ), .ZN(n3443) );
  MUX4ND0BWP U5186 ( .I0(\srf/regTable[4][6] ), .I1(\srf/regTable[5][6] ), 
        .I2(\srf/regTable[6][6] ), .I3(\srf/regTable[7][6] ), .S0(n5516), .S1(
        \srf/N16 ), .ZN(n3444) );
  MUX2ND0BWP U5187 ( .I0(n3445), .I1(n3446), .S(n5496), .ZN(\srf/N30 ) );
  MUX4ND0BWP U5188 ( .I0(\srf/regTable[0][5] ), .I1(\srf/regTable[1][5] ), 
        .I2(\srf/regTable[2][5] ), .I3(\srf/regTable[3][5] ), .S0(n5517), .S1(
        \srf/N16 ), .ZN(n3445) );
  MUX4ND0BWP U5189 ( .I0(\srf/regTable[4][5] ), .I1(\srf/regTable[5][5] ), 
        .I2(\srf/regTable[6][5] ), .I3(\srf/regTable[7][5] ), .S0(n5518), .S1(
        \srf/N16 ), .ZN(n3446) );
  MUX2ND0BWP U5190 ( .I0(n3447), .I1(n3448), .S(n5490), .ZN(\srf/N31 ) );
  MUX4ND0BWP U5191 ( .I0(\srf/regTable[0][4] ), .I1(\srf/regTable[1][4] ), 
        .I2(\srf/regTable[2][4] ), .I3(\srf/regTable[3][4] ), .S0(n5519), .S1(
        \srf/N16 ), .ZN(n3447) );
  MUX4ND0BWP U5192 ( .I0(\srf/regTable[4][4] ), .I1(\srf/regTable[5][4] ), 
        .I2(\srf/regTable[6][4] ), .I3(\srf/regTable[7][4] ), .S0(n5520), .S1(
        \srf/N16 ), .ZN(n3448) );
  MUX2ND0BWP U5193 ( .I0(n3449), .I1(n3450), .S(n5489), .ZN(\srf/N32 ) );
  MUX4ND0BWP U5194 ( .I0(\srf/regTable[0][3] ), .I1(\srf/regTable[1][3] ), 
        .I2(\srf/regTable[2][3] ), .I3(\srf/regTable[3][3] ), .S0(n5521), .S1(
        \srf/N16 ), .ZN(n3449) );
  MUX4ND0BWP U5195 ( .I0(\srf/regTable[4][3] ), .I1(\srf/regTable[5][3] ), 
        .I2(\srf/regTable[6][3] ), .I3(\srf/regTable[7][3] ), .S0(n5522), .S1(
        \srf/N16 ), .ZN(n3450) );
  MUX2ND0BWP U5196 ( .I0(n3451), .I1(n3452), .S(n5488), .ZN(\srf/N33 ) );
  MUX4ND0BWP U5197 ( .I0(\srf/regTable[0][2] ), .I1(\srf/regTable[1][2] ), 
        .I2(\srf/regTable[2][2] ), .I3(\srf/regTable[3][2] ), .S0(n5523), .S1(
        \srf/N16 ), .ZN(n3451) );
  MUX4ND0BWP U5198 ( .I0(\srf/regTable[4][2] ), .I1(\srf/regTable[5][2] ), 
        .I2(\srf/regTable[6][2] ), .I3(\srf/regTable[7][2] ), .S0(n5502), .S1(
        \srf/N16 ), .ZN(n3452) );
  MUX2ND0BWP U5199 ( .I0(n3453), .I1(n3454), .S(n5487), .ZN(\srf/N34 ) );
  MUX4ND0BWP U5200 ( .I0(\srf/regTable[0][1] ), .I1(\srf/regTable[1][1] ), 
        .I2(\srf/regTable[2][1] ), .I3(\srf/regTable[3][1] ), .S0(n5499), .S1(
        \srf/N16 ), .ZN(n3453) );
  MUX4ND0BWP U5201 ( .I0(\srf/regTable[4][1] ), .I1(\srf/regTable[5][1] ), 
        .I2(\srf/regTable[6][1] ), .I3(\srf/regTable[7][1] ), .S0(n5500), .S1(
        \srf/N16 ), .ZN(n3454) );
  MUX2ND0BWP U5202 ( .I0(n3455), .I1(n3456), .S(n5486), .ZN(\srf/N35 ) );
  MUX4ND0BWP U5203 ( .I0(\srf/regTable[0][0] ), .I1(\srf/regTable[1][0] ), 
        .I2(\srf/regTable[2][0] ), .I3(\srf/regTable[3][0] ), .S0(n5497), .S1(
        \srf/N16 ), .ZN(n3455) );
  MUX4ND0BWP U5204 ( .I0(\srf/regTable[4][0] ), .I1(\srf/regTable[5][0] ), 
        .I2(\srf/regTable[6][0] ), .I3(\srf/regTable[7][0] ), .S0(n5498), .S1(
        \srf/N16 ), .ZN(n3456) );
  MUX3ND0BWP U5205 ( .I0(\alu/N657 ), .I1(\alu/N1010 ), .I2(n5430), .S0(
        func[3]), .S1(func[0]), .ZN(n5431) );
  IND2D1BWP U5206 ( .A1(func[3]), .B1(n5475), .ZN(n5433) );
  IND2D1BWP U5207 ( .A1(func[3]), .B1(\alu/N1010 ), .ZN(n5432) );
  MUX3ND0BWP U5208 ( .I0(\alu/N658 ), .I1(\alu/N1011 ), .I2(n5434), .S0(
        func[3]), .S1(func[0]), .ZN(n5435) );
  IND2D1BWP U5209 ( .A1(func[3]), .B1(n5476), .ZN(n5437) );
  IND2D1BWP U5210 ( .A1(func[3]), .B1(\alu/N1011 ), .ZN(n5436) );
  MUX3ND0BWP U5211 ( .I0(\alu/N659 ), .I1(\alu/N1012 ), .I2(n5438), .S0(
        func[3]), .S1(func[0]), .ZN(n5439) );
  IND2D1BWP U5212 ( .A1(func[3]), .B1(n5477), .ZN(n5441) );
  IND2D1BWP U5213 ( .A1(func[3]), .B1(\alu/N1012 ), .ZN(n5440) );
  MUX3ND0BWP U5214 ( .I0(\alu/N660 ), .I1(\alu/N1013 ), .I2(n5442), .S0(
        func[3]), .S1(func[0]), .ZN(n5443) );
  IND2D1BWP U5215 ( .A1(func[3]), .B1(n5478), .ZN(n5445) );
  IND2D1BWP U5216 ( .A1(func[3]), .B1(\alu/N1013 ), .ZN(n5444) );
  MUX3ND0BWP U5217 ( .I0(\alu/N656 ), .I1(\alu/N1009 ), .I2(n5426), .S0(
        func[3]), .S1(func[0]), .ZN(n5427) );
  IND2D1BWP U5218 ( .A1(func[3]), .B1(n5474), .ZN(n5429) );
  IND2D1BWP U5219 ( .A1(func[3]), .B1(\alu/N1009 ), .ZN(n5428) );
  MUX3ND0BWP U5220 ( .I0(\alu/N655 ), .I1(\alu/N1008 ), .I2(n5422), .S0(
        func[3]), .S1(func[0]), .ZN(n5423) );
  IND2D1BWP U5221 ( .A1(func[3]), .B1(n5473), .ZN(n5425) );
  IND2D1BWP U5222 ( .A1(func[3]), .B1(\alu/N1008 ), .ZN(n5424) );
  MUX3ND0BWP U5223 ( .I0(\alu/N654 ), .I1(\alu/N1007 ), .I2(n5418), .S0(
        func[3]), .S1(func[0]), .ZN(n5419) );
  IND2D1BWP U5224 ( .A1(func[3]), .B1(n5472), .ZN(n5421) );
  IND2D1BWP U5225 ( .A1(func[3]), .B1(\alu/N1007 ), .ZN(n5420) );
  MUX3ND0BWP U5226 ( .I0(\alu/N653 ), .I1(\alu/N1006 ), .I2(n5414), .S0(
        func[3]), .S1(func[0]), .ZN(n5415) );
  IND2D1BWP U5227 ( .A1(func[3]), .B1(n5471), .ZN(n5417) );
  IND2D1BWP U5228 ( .A1(func[3]), .B1(\alu/N1006 ), .ZN(n5416) );
  MUX3ND0BWP U5229 ( .I0(\alu/N652 ), .I1(\alu/N1005 ), .I2(n5410), .S0(
        func[3]), .S1(func[0]), .ZN(n5411) );
  IND2D1BWP U5230 ( .A1(func[3]), .B1(n5470), .ZN(n5413) );
  IND2D1BWP U5231 ( .A1(func[3]), .B1(\alu/N1005 ), .ZN(n5412) );
  MUX3ND0BWP U5232 ( .I0(n3457), .I1(n5467), .I2(n3458), .S0(func[2]), .S1(
        func[1]), .ZN(result[15]) );
  MUX3ND0BWP U5233 ( .I0(\alu/N634 ), .I1(\alu/N1019 ), .I2(n5484), .S0(
        func[3]), .S1(func[0]), .ZN(n3457) );
  MUX3D1BWP U5234 ( .I0(n5466), .I1(n5467), .I2(n5468), .S0(func[0]), .S1(
        func[2]), .Z(n3458) );
  INVD1BWP U5235 ( .I(func[3]), .ZN(n5485) );
  IND2D1BWP U5236 ( .A1(func[3]), .B1(\alu/N814 ), .ZN(n5466) );
  MUX4D1BWP U5237 ( .I0(\alu/N836 ), .I1(\alu/N1018 ), .I2(\alu/N851 ), .I3(
        op2[6]), .S0(func[0]), .S1(func[2]), .Z(n5483) );
  MUX4D1BWP U5238 ( .I0(\alu/N835 ), .I1(\alu/N1017 ), .I2(op1[13]), .I3(
        op2[5]), .S0(func[0]), .S1(func[2]), .Z(n5482) );
  MUX4D1BWP U5239 ( .I0(\alu/N834 ), .I1(\alu/N1016 ), .I2(op1[12]), .I3(
        op2[4]), .S0(func[0]), .S1(func[2]), .Z(n5481) );
  MUX4D1BWP U5240 ( .I0(\alu/N833 ), .I1(\alu/N1015 ), .I2(op1[11]), .I3(
        op2[3]), .S0(func[0]), .S1(func[2]), .Z(n5480) );
  MUX4D1BWP U5241 ( .I0(\alu/N999 ), .I1(\alu/N1014 ), .I2(op1[10]), .I3(
        op2[2]), .S0(func[0]), .S1(func[2]), .Z(n5479) );
  MUX4D1BWP U5242 ( .I0(\alu/N991 ), .I1(\alu/N1013 ), .I2(op1[9]), .I3(op2[1]), .S0(func[0]), .S1(func[2]), .Z(n5478) );
  MUX4D1BWP U5243 ( .I0(\alu/N990 ), .I1(\alu/N1012 ), .I2(op1[8]), .I3(op2[0]), .S0(func[0]), .S1(func[2]), .Z(n5477) );
  MUX4D1BWP U5244 ( .I0(\alu/N989 ), .I1(\alu/N1011 ), .I2(op2[7]), .I3(op1[7]), .S0(func[0]), .S1(func[2]), .Z(n5476) );
  MUX4D1BWP U5245 ( .I0(\alu/N988 ), .I1(\alu/N1010 ), .I2(op2[6]), .I3(op1[6]), .S0(func[0]), .S1(func[2]), .Z(n5475) );
  MUX4D1BWP U5246 ( .I0(\alu/N987 ), .I1(\alu/N1009 ), .I2(op2[5]), .I3(op1[5]), .S0(func[0]), .S1(func[2]), .Z(n5474) );
  MUX4D1BWP U5247 ( .I0(\alu/N986 ), .I1(\alu/N1008 ), .I2(op2[4]), .I3(op1[4]), .S0(func[0]), .S1(func[2]), .Z(n5473) );
  MUX4D1BWP U5248 ( .I0(\alu/N985 ), .I1(\alu/N1007 ), .I2(op2[3]), .I3(op1[3]), .S0(func[0]), .S1(func[2]), .Z(n5472) );
  MUX4D1BWP U5249 ( .I0(\alu/N984 ), .I1(\alu/N1006 ), .I2(op2[2]), .I3(op1[2]), .S0(func[0]), .S1(func[2]), .Z(n5471) );
  MUX4D1BWP U5250 ( .I0(\alu/N983 ), .I1(\alu/N1005 ), .I2(op2[1]), .I3(op1[1]), .S0(func[0]), .S1(func[2]), .Z(n5470) );
  MUX4D1BWP U5251 ( .I0(\alu/N982 ), .I1(\alu/N1004 ), .I2(op2[0]), .I3(op1[0]), .S0(func[0]), .S1(func[2]), .Z(n5469) );
  IND2D1BWP U5252 ( .A1(func[3]), .B1(\alu/N1019 ), .ZN(n5467) );
  MUX3ND0BWP U5253 ( .I0(n5451), .I1(n5452), .I2(n5453), .S0(func[2]), .S1(
        func[1]), .ZN(result[11]) );
  MUX3ND0BWP U5254 ( .I0(\alu/N662 ), .I1(\alu/N1015 ), .I2(n5450), .S0(
        func[3]), .S1(func[0]), .ZN(n5451) );
  IND2D1BWP U5255 ( .A1(func[3]), .B1(n5480), .ZN(n5453) );
  IND2D1BWP U5256 ( .A1(func[3]), .B1(\alu/N1015 ), .ZN(n5452) );
  MUX3ND0BWP U5257 ( .I0(n5455), .I1(n5456), .I2(n5457), .S0(func[2]), .S1(
        func[1]), .ZN(result[12]) );
  MUX3ND0BWP U5258 ( .I0(\alu/N663 ), .I1(\alu/N1016 ), .I2(n5454), .S0(
        func[3]), .S1(func[0]), .ZN(n5455) );
  IND2D1BWP U5259 ( .A1(func[3]), .B1(n5481), .ZN(n5457) );
  IND2D1BWP U5260 ( .A1(func[3]), .B1(\alu/N1016 ), .ZN(n5456) );
  MUX3ND0BWP U5261 ( .I0(n5459), .I1(n5460), .I2(n5461), .S0(func[2]), .S1(
        func[1]), .ZN(result[13]) );
  MUX3ND0BWP U5262 ( .I0(\alu/N664 ), .I1(\alu/N1017 ), .I2(n5458), .S0(
        func[3]), .S1(func[0]), .ZN(n5459) );
  IND2D1BWP U5263 ( .A1(func[3]), .B1(n5482), .ZN(n5461) );
  IND2D1BWP U5264 ( .A1(func[3]), .B1(\alu/N1017 ), .ZN(n5460) );
  MUX3ND0BWP U5265 ( .I0(n5463), .I1(n5464), .I2(n5465), .S0(func[2]), .S1(
        func[1]), .ZN(result[14]) );
  MUX3ND0BWP U5266 ( .I0(\alu/N665 ), .I1(\alu/N1018 ), .I2(n5462), .S0(
        func[3]), .S1(func[0]), .ZN(n5463) );
  IND2D1BWP U5267 ( .A1(func[3]), .B1(n5483), .ZN(n5465) );
  IND2D1BWP U5268 ( .A1(func[3]), .B1(\alu/N1018 ), .ZN(n5464) );
  MUX3ND0BWP U5269 ( .I0(n5447), .I1(n5448), .I2(n5449), .S0(func[2]), .S1(
        func[1]), .ZN(result[10]) );
  MUX3ND0BWP U5270 ( .I0(\alu/N661 ), .I1(\alu/N1014 ), .I2(n5446), .S0(
        func[3]), .S1(func[0]), .ZN(n5447) );
  IND2D1BWP U5271 ( .A1(func[3]), .B1(n5479), .ZN(n5449) );
  IND2D1BWP U5272 ( .A1(func[3]), .B1(\alu/N1014 ), .ZN(n5448) );
  MUX3ND0BWP U5273 ( .I0(\alu/N651 ), .I1(\alu/N1004 ), .I2(n5406), .S0(
        func[3]), .S1(func[0]), .ZN(n5407) );
  IND2D1BWP U5274 ( .A1(func[3]), .B1(n5469), .ZN(n5409) );
  IND2D1BWP U5275 ( .A1(func[3]), .B1(\alu/N1004 ), .ZN(n5408) );
  MUX2D1BWP U5276 ( .I0(n3460), .I1(n3461), .S(n5070), .Z(n3459) );
  MUX4ND0BWP U5277 ( .I0(\vrf/regTable[0][35] ), .I1(\vrf/regTable[1][35] ), 
        .I2(\vrf/regTable[2][35] ), .I3(\vrf/regTable[3][35] ), .S0(n4933), 
        .S1(n5003), .ZN(n3460) );
  MUX4ND0BWP U5278 ( .I0(\vrf/regTable[4][35] ), .I1(\vrf/regTable[5][35] ), 
        .I2(\vrf/regTable[6][35] ), .I3(\vrf/regTable[7][35] ), .S0(n4933), 
        .S1(n5003), .ZN(n3461) );
  MUX2D1BWP U5279 ( .I0(n3463), .I1(n3464), .S(n5071), .Z(n3462) );
  MUX4ND0BWP U5280 ( .I0(\vrf/regTable[0][36] ), .I1(\vrf/regTable[1][36] ), 
        .I2(\vrf/regTable[2][36] ), .I3(\vrf/regTable[3][36] ), .S0(n4934), 
        .S1(n5004), .ZN(n3463) );
  MUX4ND0BWP U5281 ( .I0(\vrf/regTable[4][36] ), .I1(\vrf/regTable[5][36] ), 
        .I2(\vrf/regTable[6][36] ), .I3(\vrf/regTable[7][36] ), .S0(n4934), 
        .S1(n5004), .ZN(n3464) );
  MUX2D1BWP U5282 ( .I0(n3466), .I1(n3467), .S(n5084), .Z(n3465) );
  MUX4ND0BWP U5283 ( .I0(\vrf/regTable[0][195] ), .I1(\vrf/regTable[1][195] ), 
        .I2(\vrf/regTable[2][195] ), .I3(\vrf/regTable[3][195] ), .S0(n4960), 
        .S1(n5030), .ZN(n3466) );
  MUX4ND0BWP U5284 ( .I0(\vrf/regTable[4][195] ), .I1(\vrf/regTable[5][195] ), 
        .I2(\vrf/regTable[6][195] ), .I3(\vrf/regTable[7][195] ), .S0(n4960), 
        .S1(n5030), .ZN(n3467) );
  MUX2D1BWP U5285 ( .I0(n3469), .I1(n3470), .S(n5084), .Z(n3468) );
  MUX4ND0BWP U5286 ( .I0(\vrf/regTable[0][196] ), .I1(\vrf/regTable[1][196] ), 
        .I2(\vrf/regTable[2][196] ), .I3(\vrf/regTable[3][196] ), .S0(n4960), 
        .S1(n5030), .ZN(n3469) );
  MUX4ND0BWP U5287 ( .I0(\vrf/regTable[4][196] ), .I1(\vrf/regTable[5][196] ), 
        .I2(\vrf/regTable[6][196] ), .I3(\vrf/regTable[7][196] ), .S0(n4960), 
        .S1(n5030), .ZN(n3470) );
  MUX2D1BWP U5288 ( .I0(n3472), .I1(n3473), .S(n5082), .Z(n3471) );
  MUX4ND0BWP U5289 ( .I0(\vrf/regTable[0][176] ), .I1(\vrf/regTable[1][176] ), 
        .I2(\vrf/regTable[2][176] ), .I3(\vrf/regTable[3][176] ), .S0(n4957), 
        .S1(n5027), .ZN(n3472) );
  MUX4ND0BWP U5290 ( .I0(\vrf/regTable[4][176] ), .I1(\vrf/regTable[5][176] ), 
        .I2(\vrf/regTable[6][176] ), .I3(\vrf/regTable[7][176] ), .S0(n4957), 
        .S1(n5027), .ZN(n3473) );
  MUX2D1BWP U5291 ( .I0(n3475), .I1(n3476), .S(n5082), .Z(n3474) );
  MUX4ND0BWP U5292 ( .I0(\vrf/regTable[0][177] ), .I1(\vrf/regTable[1][177] ), 
        .I2(\vrf/regTable[2][177] ), .I3(\vrf/regTable[3][177] ), .S0(n4957), 
        .S1(n5027), .ZN(n3475) );
  MUX4ND0BWP U5293 ( .I0(\vrf/regTable[4][177] ), .I1(\vrf/regTable[5][177] ), 
        .I2(\vrf/regTable[6][177] ), .I3(\vrf/regTable[7][177] ), .S0(n4957), 
        .S1(n5027), .ZN(n3476) );
  MUX2D1BWP U5294 ( .I0(n3478), .I1(n3479), .S(n5083), .Z(n3477) );
  MUX4ND0BWP U5295 ( .I0(\vrf/regTable[0][184] ), .I1(\vrf/regTable[1][184] ), 
        .I2(\vrf/regTable[2][184] ), .I3(\vrf/regTable[3][184] ), .S0(n4958), 
        .S1(n5028), .ZN(n3478) );
  MUX4ND0BWP U5296 ( .I0(\vrf/regTable[4][184] ), .I1(\vrf/regTable[5][184] ), 
        .I2(\vrf/regTable[6][184] ), .I3(\vrf/regTable[7][184] ), .S0(n4958), 
        .S1(n5028), .ZN(n3479) );
  MUX2D1BWP U5297 ( .I0(n3481), .I1(n3482), .S(n5083), .Z(n3480) );
  MUX4ND0BWP U5298 ( .I0(\vrf/regTable[0][185] ), .I1(\vrf/regTable[1][185] ), 
        .I2(\vrf/regTable[2][185] ), .I3(\vrf/regTable[3][185] ), .S0(n4958), 
        .S1(n5028), .ZN(n3481) );
  MUX4ND0BWP U5299 ( .I0(\vrf/regTable[4][185] ), .I1(\vrf/regTable[5][185] ), 
        .I2(\vrf/regTable[6][185] ), .I3(\vrf/regTable[7][185] ), .S0(n4958), 
        .S1(n5028), .ZN(n3482) );
  MUX2D1BWP U5300 ( .I0(n3484), .I1(n3485), .S(n5083), .Z(n3483) );
  MUX4ND0BWP U5301 ( .I0(\vrf/regTable[0][186] ), .I1(\vrf/regTable[1][186] ), 
        .I2(\vrf/regTable[2][186] ), .I3(\vrf/regTable[3][186] ), .S0(n4959), 
        .S1(n5029), .ZN(n3484) );
  MUX4ND0BWP U5302 ( .I0(\vrf/regTable[4][186] ), .I1(\vrf/regTable[5][186] ), 
        .I2(\vrf/regTable[6][186] ), .I3(\vrf/regTable[7][186] ), .S0(n4959), 
        .S1(n5029), .ZN(n3485) );
  MUX2D1BWP U5303 ( .I0(n3487), .I1(n3488), .S(n5083), .Z(n3486) );
  MUX4ND0BWP U5304 ( .I0(\vrf/regTable[0][187] ), .I1(\vrf/regTable[1][187] ), 
        .I2(\vrf/regTable[2][187] ), .I3(\vrf/regTable[3][187] ), .S0(n4959), 
        .S1(n5029), .ZN(n3487) );
  MUX4ND0BWP U5305 ( .I0(\vrf/regTable[4][187] ), .I1(\vrf/regTable[5][187] ), 
        .I2(\vrf/regTable[6][187] ), .I3(\vrf/regTable[7][187] ), .S0(n4959), 
        .S1(n5029), .ZN(n3488) );
  MUX2D1BWP U5306 ( .I0(n3490), .I1(n3491), .S(n5083), .Z(n3489) );
  MUX4ND0BWP U5307 ( .I0(\vrf/regTable[0][188] ), .I1(\vrf/regTable[1][188] ), 
        .I2(\vrf/regTable[2][188] ), .I3(\vrf/regTable[3][188] ), .S0(n4959), 
        .S1(n5029), .ZN(n3490) );
  MUX4ND0BWP U5308 ( .I0(\vrf/regTable[4][188] ), .I1(\vrf/regTable[5][188] ), 
        .I2(\vrf/regTable[6][188] ), .I3(\vrf/regTable[7][188] ), .S0(n4959), 
        .S1(n5029), .ZN(n3491) );
  MUX2D1BWP U5309 ( .I0(n3493), .I1(n3494), .S(n5083), .Z(n3492) );
  MUX4ND0BWP U5310 ( .I0(\vrf/regTable[0][189] ), .I1(\vrf/regTable[1][189] ), 
        .I2(\vrf/regTable[2][189] ), .I3(\vrf/regTable[3][189] ), .S0(n4959), 
        .S1(n5029), .ZN(n3493) );
  MUX4ND0BWP U5311 ( .I0(\vrf/regTable[4][189] ), .I1(\vrf/regTable[5][189] ), 
        .I2(\vrf/regTable[6][189] ), .I3(\vrf/regTable[7][189] ), .S0(n4959), 
        .S1(n5029), .ZN(n3494) );
  MUX2D1BWP U5312 ( .I0(n3496), .I1(n3497), .S(n5083), .Z(n3495) );
  MUX4ND0BWP U5313 ( .I0(\vrf/regTable[0][190] ), .I1(\vrf/regTable[1][190] ), 
        .I2(\vrf/regTable[2][190] ), .I3(\vrf/regTable[3][190] ), .S0(n4959), 
        .S1(n5029), .ZN(n3496) );
  MUX4ND0BWP U5314 ( .I0(\vrf/regTable[4][190] ), .I1(\vrf/regTable[5][190] ), 
        .I2(\vrf/regTable[6][190] ), .I3(\vrf/regTable[7][190] ), .S0(n4959), 
        .S1(n5029), .ZN(n3497) );
  MUX2D1BWP U5315 ( .I0(n3499), .I1(n3500), .S(n5083), .Z(n3498) );
  MUX4ND0BWP U5316 ( .I0(\vrf/regTable[0][191] ), .I1(\vrf/regTable[1][191] ), 
        .I2(\vrf/regTable[2][191] ), .I3(\vrf/regTable[3][191] ), .S0(n4959), 
        .S1(n5029), .ZN(n3499) );
  MUX4ND0BWP U5317 ( .I0(\vrf/regTable[4][191] ), .I1(\vrf/regTable[5][191] ), 
        .I2(\vrf/regTable[6][191] ), .I3(\vrf/regTable[7][191] ), .S0(n4959), 
        .S1(n5029), .ZN(n3500) );
  MUX2D1BWP U5318 ( .I0(n3502), .I1(n3503), .S(n5082), .Z(n3501) );
  MUX4ND0BWP U5319 ( .I0(\vrf/regTable[0][178] ), .I1(\vrf/regTable[1][178] ), 
        .I2(\vrf/regTable[2][178] ), .I3(\vrf/regTable[3][178] ), .S0(n4957), 
        .S1(n5027), .ZN(n3502) );
  MUX4ND0BWP U5320 ( .I0(\vrf/regTable[4][178] ), .I1(\vrf/regTable[5][178] ), 
        .I2(\vrf/regTable[6][178] ), .I3(\vrf/regTable[7][178] ), .S0(n4957), 
        .S1(n5027), .ZN(n3503) );
  MUX2D1BWP U5321 ( .I0(n3505), .I1(n3506), .S(n5083), .Z(n3504) );
  MUX4ND0BWP U5322 ( .I0(\vrf/regTable[0][181] ), .I1(\vrf/regTable[1][181] ), 
        .I2(\vrf/regTable[2][181] ), .I3(\vrf/regTable[3][181] ), .S0(n4958), 
        .S1(n5028), .ZN(n3505) );
  MUX4ND0BWP U5323 ( .I0(\vrf/regTable[4][181] ), .I1(\vrf/regTable[5][181] ), 
        .I2(\vrf/regTable[6][181] ), .I3(\vrf/regTable[7][181] ), .S0(n4958), 
        .S1(n5028), .ZN(n3506) );
  MUX2D1BWP U5324 ( .I0(n3508), .I1(n3509), .S(n5083), .Z(n3507) );
  MUX4ND0BWP U5325 ( .I0(\vrf/regTable[0][182] ), .I1(\vrf/regTable[1][182] ), 
        .I2(\vrf/regTable[2][182] ), .I3(\vrf/regTable[3][182] ), .S0(n4958), 
        .S1(n5028), .ZN(n3508) );
  MUX4ND0BWP U5326 ( .I0(\vrf/regTable[4][182] ), .I1(\vrf/regTable[5][182] ), 
        .I2(\vrf/regTable[6][182] ), .I3(\vrf/regTable[7][182] ), .S0(n4958), 
        .S1(n5028), .ZN(n3509) );
  MUX2D1BWP U5327 ( .I0(n3511), .I1(n3512), .S(n5083), .Z(n3510) );
  MUX4ND0BWP U5328 ( .I0(\vrf/regTable[0][183] ), .I1(\vrf/regTable[1][183] ), 
        .I2(\vrf/regTable[2][183] ), .I3(\vrf/regTable[3][183] ), .S0(n4958), 
        .S1(n5028), .ZN(n3511) );
  MUX4ND0BWP U5329 ( .I0(\vrf/regTable[4][183] ), .I1(\vrf/regTable[5][183] ), 
        .I2(\vrf/regTable[6][183] ), .I3(\vrf/regTable[7][183] ), .S0(n4958), 
        .S1(n5028), .ZN(n3512) );
  MUX2D1BWP U5330 ( .I0(n3514), .I1(n3515), .S(n5074), .Z(n3513) );
  MUX4ND0BWP U5331 ( .I0(\vrf/regTable[0][83] ), .I1(\vrf/regTable[1][83] ), 
        .I2(\vrf/regTable[2][83] ), .I3(\vrf/regTable[3][83] ), .S0(n4941), 
        .S1(n5011), .ZN(n3514) );
  MUX4ND0BWP U5332 ( .I0(\vrf/regTable[4][83] ), .I1(\vrf/regTable[5][83] ), 
        .I2(\vrf/regTable[6][83] ), .I3(\vrf/regTable[7][83] ), .S0(n4941), 
        .S1(n5011), .ZN(n3515) );
  MUX2D1BWP U5333 ( .I0(n3517), .I1(n3518), .S(n5075), .Z(n3516) );
  MUX4ND0BWP U5334 ( .I0(\vrf/regTable[0][84] ), .I1(\vrf/regTable[1][84] ), 
        .I2(\vrf/regTable[2][84] ), .I3(\vrf/regTable[3][84] ), .S0(n4942), 
        .S1(n5012), .ZN(n3517) );
  MUX4ND0BWP U5335 ( .I0(\vrf/regTable[4][84] ), .I1(\vrf/regTable[5][84] ), 
        .I2(\vrf/regTable[6][84] ), .I3(\vrf/regTable[7][84] ), .S0(n4942), 
        .S1(n5012), .ZN(n3518) );
  MUX2D1BWP U5336 ( .I0(n3520), .I1(n3521), .S(n5077), .Z(n3519) );
  MUX4ND0BWP U5337 ( .I0(\vrf/regTable[0][112] ), .I1(\vrf/regTable[1][112] ), 
        .I2(\vrf/regTable[2][112] ), .I3(\vrf/regTable[3][112] ), .S0(n4946), 
        .S1(n5016), .ZN(n3520) );
  MUX4ND0BWP U5338 ( .I0(\vrf/regTable[4][112] ), .I1(\vrf/regTable[5][112] ), 
        .I2(\vrf/regTable[6][112] ), .I3(\vrf/regTable[7][112] ), .S0(n4946), 
        .S1(n5016), .ZN(n3521) );
  MUX2D1BWP U5339 ( .I0(n3523), .I1(n3524), .S(n5077), .Z(n3522) );
  MUX4ND0BWP U5340 ( .I0(\vrf/regTable[0][113] ), .I1(\vrf/regTable[1][113] ), 
        .I2(\vrf/regTable[2][113] ), .I3(\vrf/regTable[3][113] ), .S0(n4946), 
        .S1(n5016), .ZN(n3523) );
  MUX4ND0BWP U5341 ( .I0(\vrf/regTable[4][113] ), .I1(\vrf/regTable[5][113] ), 
        .I2(\vrf/regTable[6][113] ), .I3(\vrf/regTable[7][113] ), .S0(n4946), 
        .S1(n5016), .ZN(n3524) );
  MUX2D1BWP U5342 ( .I0(n3526), .I1(n3527), .S(n5078), .Z(n3525) );
  MUX4ND0BWP U5343 ( .I0(\vrf/regTable[0][120] ), .I1(\vrf/regTable[1][120] ), 
        .I2(\vrf/regTable[2][120] ), .I3(\vrf/regTable[3][120] ), .S0(n4948), 
        .S1(n5018), .ZN(n3526) );
  MUX4ND0BWP U5344 ( .I0(\vrf/regTable[4][120] ), .I1(\vrf/regTable[5][120] ), 
        .I2(\vrf/regTable[6][120] ), .I3(\vrf/regTable[7][120] ), .S0(n4948), 
        .S1(n5018), .ZN(n3527) );
  MUX2D1BWP U5345 ( .I0(n3529), .I1(n3530), .S(n5078), .Z(n3528) );
  MUX4ND0BWP U5346 ( .I0(\vrf/regTable[0][121] ), .I1(\vrf/regTable[1][121] ), 
        .I2(\vrf/regTable[2][121] ), .I3(\vrf/regTable[3][121] ), .S0(n4948), 
        .S1(n5018), .ZN(n3529) );
  MUX4ND0BWP U5347 ( .I0(\vrf/regTable[4][121] ), .I1(\vrf/regTable[5][121] ), 
        .I2(\vrf/regTable[6][121] ), .I3(\vrf/regTable[7][121] ), .S0(n4948), 
        .S1(n5018), .ZN(n3530) );
  MUX2D1BWP U5348 ( .I0(n3532), .I1(n3533), .S(n5078), .Z(n3531) );
  MUX4ND0BWP U5349 ( .I0(\vrf/regTable[0][122] ), .I1(\vrf/regTable[1][122] ), 
        .I2(\vrf/regTable[2][122] ), .I3(\vrf/regTable[3][122] ), .S0(n4948), 
        .S1(n5018), .ZN(n3532) );
  MUX4ND0BWP U5350 ( .I0(\vrf/regTable[4][122] ), .I1(\vrf/regTable[5][122] ), 
        .I2(\vrf/regTable[6][122] ), .I3(\vrf/regTable[7][122] ), .S0(n4948), 
        .S1(n5018), .ZN(n3533) );
  MUX2D1BWP U5351 ( .I0(n3535), .I1(n3536), .S(n5078), .Z(n3534) );
  MUX4ND0BWP U5352 ( .I0(\vrf/regTable[0][123] ), .I1(\vrf/regTable[1][123] ), 
        .I2(\vrf/regTable[2][123] ), .I3(\vrf/regTable[3][123] ), .S0(n4948), 
        .S1(n5018), .ZN(n3535) );
  MUX4ND0BWP U5353 ( .I0(\vrf/regTable[4][123] ), .I1(\vrf/regTable[5][123] ), 
        .I2(\vrf/regTable[6][123] ), .I3(\vrf/regTable[7][123] ), .S0(n4948), 
        .S1(n5018), .ZN(n3536) );
  MUX2D1BWP U5354 ( .I0(n3538), .I1(n3539), .S(n5078), .Z(n3537) );
  MUX4ND0BWP U5355 ( .I0(\vrf/regTable[0][124] ), .I1(\vrf/regTable[1][124] ), 
        .I2(\vrf/regTable[2][124] ), .I3(\vrf/regTable[3][124] ), .S0(n4948), 
        .S1(n5018), .ZN(n3538) );
  MUX4ND0BWP U5356 ( .I0(\vrf/regTable[4][124] ), .I1(\vrf/regTable[5][124] ), 
        .I2(\vrf/regTable[6][124] ), .I3(\vrf/regTable[7][124] ), .S0(n4948), 
        .S1(n5018), .ZN(n3539) );
  MUX2D1BWP U5357 ( .I0(n3541), .I1(n3542), .S(n5078), .Z(n3540) );
  MUX4ND0BWP U5358 ( .I0(\vrf/regTable[0][125] ), .I1(\vrf/regTable[1][125] ), 
        .I2(\vrf/regTable[2][125] ), .I3(\vrf/regTable[3][125] ), .S0(n4948), 
        .S1(n5018), .ZN(n3541) );
  MUX4ND0BWP U5359 ( .I0(\vrf/regTable[4][125] ), .I1(\vrf/regTable[5][125] ), 
        .I2(\vrf/regTable[6][125] ), .I3(\vrf/regTable[7][125] ), .S0(n4948), 
        .S1(n5018), .ZN(n3542) );
  MUX2D1BWP U5360 ( .I0(n3544), .I1(n3545), .S(n5078), .Z(n3543) );
  MUX4ND0BWP U5361 ( .I0(\vrf/regTable[0][126] ), .I1(\vrf/regTable[1][126] ), 
        .I2(\vrf/regTable[2][126] ), .I3(\vrf/regTable[3][126] ), .S0(n4949), 
        .S1(n5019), .ZN(n3544) );
  MUX4ND0BWP U5362 ( .I0(\vrf/regTable[4][126] ), .I1(\vrf/regTable[5][126] ), 
        .I2(\vrf/regTable[6][126] ), .I3(\vrf/regTable[7][126] ), .S0(n4949), 
        .S1(n5019), .ZN(n3545) );
  MUX2D1BWP U5363 ( .I0(n3547), .I1(n3548), .S(n5078), .Z(n3546) );
  MUX4ND0BWP U5364 ( .I0(\vrf/regTable[0][127] ), .I1(\vrf/regTable[1][127] ), 
        .I2(\vrf/regTable[2][127] ), .I3(\vrf/regTable[3][127] ), .S0(n4949), 
        .S1(n5019), .ZN(n3547) );
  MUX4ND0BWP U5365 ( .I0(\vrf/regTable[4][127] ), .I1(\vrf/regTable[5][127] ), 
        .I2(\vrf/regTable[6][127] ), .I3(\vrf/regTable[7][127] ), .S0(n4949), 
        .S1(n5019), .ZN(n3548) );
  MUX2D1BWP U5366 ( .I0(n3550), .I1(n3551), .S(n5077), .Z(n3549) );
  MUX4ND0BWP U5367 ( .I0(\vrf/regTable[0][114] ), .I1(\vrf/regTable[1][114] ), 
        .I2(\vrf/regTable[2][114] ), .I3(\vrf/regTable[3][114] ), .S0(n4947), 
        .S1(n5017), .ZN(n3550) );
  MUX4ND0BWP U5368 ( .I0(\vrf/regTable[4][114] ), .I1(\vrf/regTable[5][114] ), 
        .I2(\vrf/regTable[6][114] ), .I3(\vrf/regTable[7][114] ), .S0(n4947), 
        .S1(n5017), .ZN(n3551) );
  MUX2D1BWP U5369 ( .I0(n3553), .I1(n3554), .S(n5077), .Z(n3552) );
  MUX4ND0BWP U5370 ( .I0(\vrf/regTable[0][117] ), .I1(\vrf/regTable[1][117] ), 
        .I2(\vrf/regTable[2][117] ), .I3(\vrf/regTable[3][117] ), .S0(n4947), 
        .S1(n5017), .ZN(n3553) );
  MUX4ND0BWP U5371 ( .I0(\vrf/regTable[4][117] ), .I1(\vrf/regTable[5][117] ), 
        .I2(\vrf/regTable[6][117] ), .I3(\vrf/regTable[7][117] ), .S0(n4947), 
        .S1(n5017), .ZN(n3554) );
  MUX2D1BWP U5372 ( .I0(n3556), .I1(n3557), .S(n5077), .Z(n3555) );
  MUX4ND0BWP U5373 ( .I0(\vrf/regTable[0][118] ), .I1(\vrf/regTable[1][118] ), 
        .I2(\vrf/regTable[2][118] ), .I3(\vrf/regTable[3][118] ), .S0(n4947), 
        .S1(n5017), .ZN(n3556) );
  MUX4ND0BWP U5374 ( .I0(\vrf/regTable[4][118] ), .I1(\vrf/regTable[5][118] ), 
        .I2(\vrf/regTable[6][118] ), .I3(\vrf/regTable[7][118] ), .S0(n4947), 
        .S1(n5017), .ZN(n3557) );
  MUX2D1BWP U5375 ( .I0(n3559), .I1(n3560), .S(n5077), .Z(n3558) );
  MUX4ND0BWP U5376 ( .I0(\vrf/regTable[0][119] ), .I1(\vrf/regTable[1][119] ), 
        .I2(\vrf/regTable[2][119] ), .I3(\vrf/regTable[3][119] ), .S0(n4947), 
        .S1(n5017), .ZN(n3559) );
  MUX4ND0BWP U5377 ( .I0(\vrf/regTable[4][119] ), .I1(\vrf/regTable[5][119] ), 
        .I2(\vrf/regTable[6][119] ), .I3(\vrf/regTable[7][119] ), .S0(n4947), 
        .S1(n5017), .ZN(n3560) );
  MUX2D1BWP U5378 ( .I0(n3562), .I1(n3563), .S(n5085), .Z(n3561) );
  MUX4ND0BWP U5379 ( .I0(\vrf/regTable[0][211] ), .I1(\vrf/regTable[1][211] ), 
        .I2(\vrf/regTable[2][211] ), .I3(\vrf/regTable[3][211] ), .S0(n4963), 
        .S1(n5033), .ZN(n3562) );
  MUX4ND0BWP U5380 ( .I0(\vrf/regTable[4][211] ), .I1(\vrf/regTable[5][211] ), 
        .I2(\vrf/regTable[6][211] ), .I3(\vrf/regTable[7][211] ), .S0(n4963), 
        .S1(n5033), .ZN(n3563) );
  MUX2D1BWP U5381 ( .I0(n3565), .I1(n3566), .S(n5085), .Z(n3564) );
  MUX4ND0BWP U5382 ( .I0(\vrf/regTable[0][212] ), .I1(\vrf/regTable[1][212] ), 
        .I2(\vrf/regTable[2][212] ), .I3(\vrf/regTable[3][212] ), .S0(n4963), 
        .S1(n5033), .ZN(n3565) );
  MUX4ND0BWP U5383 ( .I0(\vrf/regTable[4][212] ), .I1(\vrf/regTable[5][212] ), 
        .I2(\vrf/regTable[6][212] ), .I3(\vrf/regTable[7][212] ), .S0(n4963), 
        .S1(n5033), .ZN(n3566) );
  MUX2D1BWP U5384 ( .I0(n3568), .I1(n3569), .S(n5072), .Z(n3567) );
  MUX4ND0BWP U5385 ( .I0(\vrf/regTable[0][51] ), .I1(\vrf/regTable[1][51] ), 
        .I2(\vrf/regTable[2][51] ), .I3(\vrf/regTable[3][51] ), .S0(n4936), 
        .S1(n5006), .ZN(n3568) );
  MUX4ND0BWP U5386 ( .I0(\vrf/regTable[4][51] ), .I1(\vrf/regTable[5][51] ), 
        .I2(\vrf/regTable[6][51] ), .I3(\vrf/regTable[7][51] ), .S0(n4936), 
        .S1(n5006), .ZN(n3569) );
  MUX2D1BWP U5387 ( .I0(n3571), .I1(n3572), .S(n5072), .Z(n3570) );
  MUX4ND0BWP U5388 ( .I0(\vrf/regTable[0][52] ), .I1(\vrf/regTable[1][52] ), 
        .I2(\vrf/regTable[2][52] ), .I3(\vrf/regTable[3][52] ), .S0(n4936), 
        .S1(n5006), .ZN(n3571) );
  MUX4ND0BWP U5389 ( .I0(\vrf/regTable[4][52] ), .I1(\vrf/regTable[5][52] ), 
        .I2(\vrf/regTable[6][52] ), .I3(\vrf/regTable[7][52] ), .S0(n4936), 
        .S1(n5006), .ZN(n3572) );
  MUX2D1BWP U5390 ( .I0(n3574), .I1(n3575), .S(n5069), .Z(n3573) );
  MUX4ND0BWP U5391 ( .I0(\vrf/regTable[0][16] ), .I1(\vrf/regTable[1][16] ), 
        .I2(\vrf/regTable[2][16] ), .I3(\vrf/regTable[3][16] ), .S0(n4930), 
        .S1(n5000), .ZN(n3574) );
  MUX4ND0BWP U5392 ( .I0(\vrf/regTable[4][16] ), .I1(\vrf/regTable[5][16] ), 
        .I2(\vrf/regTable[6][16] ), .I3(\vrf/regTable[7][16] ), .S0(n4930), 
        .S1(n5000), .ZN(n3575) );
  MUX2D1BWP U5393 ( .I0(n3577), .I1(n3578), .S(n5069), .Z(n3576) );
  MUX4ND0BWP U5394 ( .I0(\vrf/regTable[0][17] ), .I1(\vrf/regTable[1][17] ), 
        .I2(\vrf/regTable[2][17] ), .I3(\vrf/regTable[3][17] ), .S0(n4930), 
        .S1(n5000), .ZN(n3577) );
  MUX4ND0BWP U5395 ( .I0(\vrf/regTable[4][17] ), .I1(\vrf/regTable[5][17] ), 
        .I2(\vrf/regTable[6][17] ), .I3(\vrf/regTable[7][17] ), .S0(n4930), 
        .S1(n5000), .ZN(n3578) );
  MUX2D1BWP U5396 ( .I0(n3580), .I1(n3581), .S(n5070), .Z(n3579) );
  MUX4ND0BWP U5397 ( .I0(\vrf/regTable[0][24] ), .I1(\vrf/regTable[1][24] ), 
        .I2(\vrf/regTable[2][24] ), .I3(\vrf/regTable[3][24] ), .S0(n4932), 
        .S1(n5002), .ZN(n3580) );
  MUX4ND0BWP U5398 ( .I0(\vrf/regTable[4][24] ), .I1(\vrf/regTable[5][24] ), 
        .I2(\vrf/regTable[6][24] ), .I3(\vrf/regTable[7][24] ), .S0(n4932), 
        .S1(n5002), .ZN(n3581) );
  MUX2D1BWP U5399 ( .I0(n3583), .I1(n3584), .S(n5070), .Z(n3582) );
  MUX4ND0BWP U5400 ( .I0(\vrf/regTable[0][25] ), .I1(\vrf/regTable[1][25] ), 
        .I2(\vrf/regTable[2][25] ), .I3(\vrf/regTable[3][25] ), .S0(n4932), 
        .S1(n5002), .ZN(n3583) );
  MUX4ND0BWP U5401 ( .I0(\vrf/regTable[4][25] ), .I1(\vrf/regTable[5][25] ), 
        .I2(\vrf/regTable[6][25] ), .I3(\vrf/regTable[7][25] ), .S0(n4932), 
        .S1(n5002), .ZN(n3584) );
  MUX2D1BWP U5402 ( .I0(n3586), .I1(n3587), .S(n5070), .Z(n3585) );
  MUX4ND0BWP U5403 ( .I0(\vrf/regTable[0][26] ), .I1(\vrf/regTable[1][26] ), 
        .I2(\vrf/regTable[2][26] ), .I3(\vrf/regTable[3][26] ), .S0(n4932), 
        .S1(n5002), .ZN(n3586) );
  MUX4ND0BWP U5404 ( .I0(\vrf/regTable[4][26] ), .I1(\vrf/regTable[5][26] ), 
        .I2(\vrf/regTable[6][26] ), .I3(\vrf/regTable[7][26] ), .S0(n4932), 
        .S1(n5002), .ZN(n3587) );
  MUX2D1BWP U5405 ( .I0(n3589), .I1(n3590), .S(n5070), .Z(n3588) );
  MUX4ND0BWP U5406 ( .I0(\vrf/regTable[0][27] ), .I1(\vrf/regTable[1][27] ), 
        .I2(\vrf/regTable[2][27] ), .I3(\vrf/regTable[3][27] ), .S0(n4932), 
        .S1(n5002), .ZN(n3589) );
  MUX4ND0BWP U5407 ( .I0(\vrf/regTable[4][27] ), .I1(\vrf/regTable[5][27] ), 
        .I2(\vrf/regTable[6][27] ), .I3(\vrf/regTable[7][27] ), .S0(n4932), 
        .S1(n5002), .ZN(n3590) );
  MUX2D1BWP U5408 ( .I0(n3592), .I1(n3593), .S(n5070), .Z(n3591) );
  MUX4ND0BWP U5409 ( .I0(\vrf/regTable[0][28] ), .I1(\vrf/regTable[1][28] ), 
        .I2(\vrf/regTable[2][28] ), .I3(\vrf/regTable[3][28] ), .S0(n4932), 
        .S1(n5002), .ZN(n3592) );
  MUX4ND0BWP U5410 ( .I0(\vrf/regTable[4][28] ), .I1(\vrf/regTable[5][28] ), 
        .I2(\vrf/regTable[6][28] ), .I3(\vrf/regTable[7][28] ), .S0(n4932), 
        .S1(n5002), .ZN(n3593) );
  MUX2D1BWP U5411 ( .I0(n3595), .I1(n3596), .S(n5070), .Z(n3594) );
  MUX4ND0BWP U5412 ( .I0(\vrf/regTable[0][29] ), .I1(\vrf/regTable[1][29] ), 
        .I2(\vrf/regTable[2][29] ), .I3(\vrf/regTable[3][29] ), .S0(n4932), 
        .S1(n5002), .ZN(n3595) );
  MUX4ND0BWP U5413 ( .I0(\vrf/regTable[4][29] ), .I1(\vrf/regTable[5][29] ), 
        .I2(\vrf/regTable[6][29] ), .I3(\vrf/regTable[7][29] ), .S0(n4932), 
        .S1(n5002), .ZN(n3596) );
  MUX2D1BWP U5414 ( .I0(n3598), .I1(n3599), .S(n5070), .Z(n3597) );
  MUX4ND0BWP U5415 ( .I0(\vrf/regTable[0][30] ), .I1(\vrf/regTable[1][30] ), 
        .I2(\vrf/regTable[2][30] ), .I3(\vrf/regTable[3][30] ), .S0(n4933), 
        .S1(n5003), .ZN(n3598) );
  MUX4ND0BWP U5416 ( .I0(\vrf/regTable[4][30] ), .I1(\vrf/regTable[5][30] ), 
        .I2(\vrf/regTable[6][30] ), .I3(\vrf/regTable[7][30] ), .S0(n4933), 
        .S1(n5003), .ZN(n3599) );
  MUX2D1BWP U5417 ( .I0(n3601), .I1(n3602), .S(n5070), .Z(n3600) );
  MUX4ND0BWP U5418 ( .I0(\vrf/regTable[0][31] ), .I1(\vrf/regTable[1][31] ), 
        .I2(\vrf/regTable[2][31] ), .I3(\vrf/regTable[3][31] ), .S0(n4933), 
        .S1(n5003), .ZN(n3601) );
  MUX4ND0BWP U5419 ( .I0(\vrf/regTable[4][31] ), .I1(\vrf/regTable[5][31] ), 
        .I2(\vrf/regTable[6][31] ), .I3(\vrf/regTable[7][31] ), .S0(n4933), 
        .S1(n5003), .ZN(n3602) );
  MUX2D1BWP U5420 ( .I0(n3604), .I1(n3605), .S(n5069), .Z(n3603) );
  MUX4ND0BWP U5421 ( .I0(\vrf/regTable[0][18] ), .I1(\vrf/regTable[1][18] ), 
        .I2(\vrf/regTable[2][18] ), .I3(\vrf/regTable[3][18] ), .S0(n4931), 
        .S1(n5001), .ZN(n3604) );
  MUX4ND0BWP U5422 ( .I0(\vrf/regTable[4][18] ), .I1(\vrf/regTable[5][18] ), 
        .I2(\vrf/regTable[6][18] ), .I3(\vrf/regTable[7][18] ), .S0(n4931), 
        .S1(n5001), .ZN(n3605) );
  MUX2D1BWP U5423 ( .I0(n3607), .I1(n3608), .S(n5069), .Z(n3606) );
  MUX4ND0BWP U5424 ( .I0(\vrf/regTable[0][21] ), .I1(\vrf/regTable[1][21] ), 
        .I2(\vrf/regTable[2][21] ), .I3(\vrf/regTable[3][21] ), .S0(n4931), 
        .S1(n5001), .ZN(n3607) );
  MUX4ND0BWP U5425 ( .I0(\vrf/regTable[4][21] ), .I1(\vrf/regTable[5][21] ), 
        .I2(\vrf/regTable[6][21] ), .I3(\vrf/regTable[7][21] ), .S0(n4931), 
        .S1(n5001), .ZN(n3608) );
  MUX2D1BWP U5426 ( .I0(n3610), .I1(n3611), .S(n5069), .Z(n3609) );
  MUX4ND0BWP U5427 ( .I0(\vrf/regTable[0][22] ), .I1(\vrf/regTable[1][22] ), 
        .I2(\vrf/regTable[2][22] ), .I3(\vrf/regTable[3][22] ), .S0(n4931), 
        .S1(n5001), .ZN(n3610) );
  MUX4ND0BWP U5428 ( .I0(\vrf/regTable[4][22] ), .I1(\vrf/regTable[5][22] ), 
        .I2(\vrf/regTable[6][22] ), .I3(\vrf/regTable[7][22] ), .S0(n4931), 
        .S1(n5001), .ZN(n3611) );
  MUX2D1BWP U5429 ( .I0(n3613), .I1(n3614), .S(n5069), .Z(n3612) );
  MUX4ND0BWP U5430 ( .I0(\vrf/regTable[0][23] ), .I1(\vrf/regTable[1][23] ), 
        .I2(\vrf/regTable[2][23] ), .I3(\vrf/regTable[3][23] ), .S0(n4931), 
        .S1(n5001), .ZN(n3613) );
  MUX4ND0BWP U5431 ( .I0(\vrf/regTable[4][23] ), .I1(\vrf/regTable[5][23] ), 
        .I2(\vrf/regTable[6][23] ), .I3(\vrf/regTable[7][23] ), .S0(n4931), 
        .S1(n5001), .ZN(n3614) );
  MUX2D1BWP U5432 ( .I0(n3616), .I1(n3617), .S(n5076), .Z(n3615) );
  MUX4ND0BWP U5433 ( .I0(\vrf/regTable[0][99] ), .I1(\vrf/regTable[1][99] ), 
        .I2(\vrf/regTable[2][99] ), .I3(\vrf/regTable[3][99] ), .S0(n4944), 
        .S1(n5014), .ZN(n3616) );
  MUX4ND0BWP U5434 ( .I0(\vrf/regTable[4][99] ), .I1(\vrf/regTable[5][99] ), 
        .I2(\vrf/regTable[6][99] ), .I3(\vrf/regTable[7][99] ), .S0(n4944), 
        .S1(n5014), .ZN(n3617) );
  MUX2D1BWP U5435 ( .I0(n3619), .I1(n3620), .S(n5076), .Z(n3618) );
  MUX4ND0BWP U5436 ( .I0(\vrf/regTable[0][100] ), .I1(\vrf/regTable[1][100] ), 
        .I2(\vrf/regTable[2][100] ), .I3(\vrf/regTable[3][100] ), .S0(n4944), 
        .S1(n5014), .ZN(n3619) );
  MUX4ND0BWP U5437 ( .I0(\vrf/regTable[4][100] ), .I1(\vrf/regTable[5][100] ), 
        .I2(\vrf/regTable[6][100] ), .I3(\vrf/regTable[7][100] ), .S0(n4944), 
        .S1(n5014), .ZN(n3620) );
  MUX2D1BWP U5438 ( .I0(n3622), .I1(n3623), .S(n5073), .Z(n3621) );
  MUX4ND0BWP U5439 ( .I0(\vrf/regTable[0][67] ), .I1(\vrf/regTable[1][67] ), 
        .I2(\vrf/regTable[2][67] ), .I3(\vrf/regTable[3][67] ), .S0(n4939), 
        .S1(n5009), .ZN(n3622) );
  MUX4ND0BWP U5440 ( .I0(\vrf/regTable[4][67] ), .I1(\vrf/regTable[5][67] ), 
        .I2(\vrf/regTable[6][67] ), .I3(\vrf/regTable[7][67] ), .S0(n4939), 
        .S1(n5009), .ZN(n3623) );
  MUX2D1BWP U5441 ( .I0(n3625), .I1(n3626), .S(n5073), .Z(n3624) );
  MUX4ND0BWP U5442 ( .I0(\vrf/regTable[0][68] ), .I1(\vrf/regTable[1][68] ), 
        .I2(\vrf/regTable[2][68] ), .I3(\vrf/regTable[3][68] ), .S0(n4939), 
        .S1(n5009), .ZN(n3625) );
  MUX4ND0BWP U5443 ( .I0(\vrf/regTable[4][68] ), .I1(\vrf/regTable[5][68] ), 
        .I2(\vrf/regTable[6][68] ), .I3(\vrf/regTable[7][68] ), .S0(n4939), 
        .S1(n5009), .ZN(n3626) );
  MUX2D1BWP U5444 ( .I0(n3628), .I1(n3629), .S(n5081), .Z(n3627) );
  MUX4ND0BWP U5445 ( .I0(\vrf/regTable[0][163] ), .I1(\vrf/regTable[1][163] ), 
        .I2(\vrf/regTable[2][163] ), .I3(\vrf/regTable[3][163] ), .S0(n4955), 
        .S1(n5025), .ZN(n3628) );
  MUX4ND0BWP U5446 ( .I0(\vrf/regTable[4][163] ), .I1(\vrf/regTable[5][163] ), 
        .I2(\vrf/regTable[6][163] ), .I3(\vrf/regTable[7][163] ), .S0(n4955), 
        .S1(n5025), .ZN(n3629) );
  MUX2D1BWP U5447 ( .I0(n3631), .I1(n3632), .S(n5081), .Z(n3630) );
  MUX4ND0BWP U5448 ( .I0(\vrf/regTable[0][164] ), .I1(\vrf/regTable[1][164] ), 
        .I2(\vrf/regTable[2][164] ), .I3(\vrf/regTable[3][164] ), .S0(n4955), 
        .S1(n5025), .ZN(n3631) );
  MUX4ND0BWP U5449 ( .I0(\vrf/regTable[4][164] ), .I1(\vrf/regTable[5][164] ), 
        .I2(\vrf/regTable[6][164] ), .I3(\vrf/regTable[7][164] ), .S0(n4955), 
        .S1(n5025), .ZN(n3632) );
  MUX2D1BWP U5450 ( .I0(n3634), .I1(n3635), .S(n5068), .Z(n3633) );
  MUX4ND0BWP U5451 ( .I0(\vrf/regTable[0][11] ), .I1(\vrf/regTable[1][11] ), 
        .I2(\vrf/regTable[2][11] ), .I3(\vrf/regTable[3][11] ), .S0(n4929), 
        .S1(n4999), .ZN(n3634) );
  MUX4ND0BWP U5452 ( .I0(\vrf/regTable[4][11] ), .I1(\vrf/regTable[5][11] ), 
        .I2(\vrf/regTable[6][11] ), .I3(\vrf/regTable[7][11] ), .S0(n4929), 
        .S1(n4999), .ZN(n3635) );
  MUX2D1BWP U5453 ( .I0(n3637), .I1(n3638), .S(n5069), .Z(n3636) );
  MUX4ND0BWP U5454 ( .I0(\vrf/regTable[0][12] ), .I1(\vrf/regTable[1][12] ), 
        .I2(\vrf/regTable[2][12] ), .I3(\vrf/regTable[3][12] ), .S0(n4930), 
        .S1(n5000), .ZN(n3637) );
  MUX4ND0BWP U5455 ( .I0(\vrf/regTable[4][12] ), .I1(\vrf/regTable[5][12] ), 
        .I2(\vrf/regTable[6][12] ), .I3(\vrf/regTable[7][12] ), .S0(n4930), 
        .S1(n5000), .ZN(n3638) );
  MUX2D1BWP U5456 ( .I0(n3640), .I1(n3641), .S(n5069), .Z(n3639) );
  MUX4ND0BWP U5457 ( .I0(\vrf/regTable[0][13] ), .I1(\vrf/regTable[1][13] ), 
        .I2(\vrf/regTable[2][13] ), .I3(\vrf/regTable[3][13] ), .S0(n4930), 
        .S1(n5000), .ZN(n3640) );
  MUX4ND0BWP U5458 ( .I0(\vrf/regTable[4][13] ), .I1(\vrf/regTable[5][13] ), 
        .I2(\vrf/regTable[6][13] ), .I3(\vrf/regTable[7][13] ), .S0(n4930), 
        .S1(n5000), .ZN(n3641) );
  MUX2D1BWP U5459 ( .I0(n3643), .I1(n3644), .S(n5069), .Z(n3642) );
  MUX4ND0BWP U5460 ( .I0(\vrf/regTable[0][14] ), .I1(\vrf/regTable[1][14] ), 
        .I2(\vrf/regTable[2][14] ), .I3(\vrf/regTable[3][14] ), .S0(n4930), 
        .S1(n5000), .ZN(n3643) );
  MUX4ND0BWP U5461 ( .I0(\vrf/regTable[4][14] ), .I1(\vrf/regTable[5][14] ), 
        .I2(\vrf/regTable[6][14] ), .I3(\vrf/regTable[7][14] ), .S0(n4930), 
        .S1(n5000), .ZN(n3644) );
  MUX2D1BWP U5462 ( .I0(n3646), .I1(n3647), .S(n5069), .Z(n3645) );
  MUX4ND0BWP U5463 ( .I0(\vrf/regTable[0][15] ), .I1(\vrf/regTable[1][15] ), 
        .I2(\vrf/regTable[2][15] ), .I3(\vrf/regTable[3][15] ), .S0(n4930), 
        .S1(n5000), .ZN(n3646) );
  MUX4ND0BWP U5464 ( .I0(\vrf/regTable[4][15] ), .I1(\vrf/regTable[5][15] ), 
        .I2(\vrf/regTable[6][15] ), .I3(\vrf/regTable[7][15] ), .S0(n4930), 
        .S1(n5000), .ZN(n3647) );
  MUX2D1BWP U5465 ( .I0(n3649), .I1(n3650), .S(n5068), .Z(n3648) );
  MUX4ND0BWP U5466 ( .I0(\vrf/regTable[0][0] ), .I1(\vrf/regTable[1][0] ), 
        .I2(\vrf/regTable[2][0] ), .I3(\vrf/regTable[3][0] ), .S0(n4928), .S1(
        n4998), .ZN(n3649) );
  MUX4ND0BWP U5467 ( .I0(\vrf/regTable[4][0] ), .I1(\vrf/regTable[5][0] ), 
        .I2(\vrf/regTable[6][0] ), .I3(\vrf/regTable[7][0] ), .S0(n4928), .S1(
        n4998), .ZN(n3650) );
  MUX2D1BWP U5468 ( .I0(n3652), .I1(n3653), .S(n5068), .Z(n3651) );
  MUX4ND0BWP U5469 ( .I0(\vrf/regTable[0][1] ), .I1(\vrf/regTable[1][1] ), 
        .I2(\vrf/regTable[2][1] ), .I3(\vrf/regTable[3][1] ), .S0(n4928), .S1(
        n4998), .ZN(n3652) );
  MUX4ND0BWP U5470 ( .I0(\vrf/regTable[4][1] ), .I1(\vrf/regTable[5][1] ), 
        .I2(\vrf/regTable[6][1] ), .I3(\vrf/regTable[7][1] ), .S0(n4928), .S1(
        n4998), .ZN(n3653) );
  MUX2D1BWP U5471 ( .I0(n3655), .I1(n3656), .S(n5068), .Z(n3654) );
  MUX4ND0BWP U5472 ( .I0(\vrf/regTable[0][2] ), .I1(\vrf/regTable[1][2] ), 
        .I2(\vrf/regTable[2][2] ), .I3(\vrf/regTable[3][2] ), .S0(n4928), .S1(
        n4998), .ZN(n3655) );
  MUX4ND0BWP U5473 ( .I0(\vrf/regTable[4][2] ), .I1(\vrf/regTable[5][2] ), 
        .I2(\vrf/regTable[6][2] ), .I3(\vrf/regTable[7][2] ), .S0(n4928), .S1(
        n4998), .ZN(n3656) );
  MUX2D1BWP U5474 ( .I0(n3658), .I1(n3659), .S(n5068), .Z(n3657) );
  MUX4ND0BWP U5475 ( .I0(\vrf/regTable[0][5] ), .I1(\vrf/regTable[1][5] ), 
        .I2(\vrf/regTable[2][5] ), .I3(\vrf/regTable[3][5] ), .S0(n4928), .S1(
        n4998), .ZN(n3658) );
  MUX4ND0BWP U5476 ( .I0(\vrf/regTable[4][5] ), .I1(\vrf/regTable[5][5] ), 
        .I2(\vrf/regTable[6][5] ), .I3(\vrf/regTable[7][5] ), .S0(n4928), .S1(
        n4998), .ZN(n3659) );
  MUX2D1BWP U5477 ( .I0(n3661), .I1(n3662), .S(n5068), .Z(n3660) );
  MUX4ND0BWP U5478 ( .I0(\vrf/regTable[0][6] ), .I1(\vrf/regTable[1][6] ), 
        .I2(\vrf/regTable[2][6] ), .I3(\vrf/regTable[3][6] ), .S0(n4929), .S1(
        n4999), .ZN(n3661) );
  MUX4ND0BWP U5479 ( .I0(\vrf/regTable[4][6] ), .I1(\vrf/regTable[5][6] ), 
        .I2(\vrf/regTable[6][6] ), .I3(\vrf/regTable[7][6] ), .S0(n4929), .S1(
        n4999), .ZN(n3662) );
  MUX2D1BWP U5480 ( .I0(n3664), .I1(n3665), .S(n5068), .Z(n3663) );
  MUX4ND0BWP U5481 ( .I0(\vrf/regTable[0][7] ), .I1(\vrf/regTable[1][7] ), 
        .I2(\vrf/regTable[2][7] ), .I3(\vrf/regTable[3][7] ), .S0(n4929), .S1(
        n4999), .ZN(n3664) );
  MUX4ND0BWP U5482 ( .I0(\vrf/regTable[4][7] ), .I1(\vrf/regTable[5][7] ), 
        .I2(\vrf/regTable[6][7] ), .I3(\vrf/regTable[7][7] ), .S0(n4929), .S1(
        n4999), .ZN(n3665) );
  MUX2D1BWP U5483 ( .I0(n3667), .I1(n3668), .S(n5068), .Z(n3666) );
  MUX4ND0BWP U5484 ( .I0(\vrf/regTable[0][8] ), .I1(\vrf/regTable[1][8] ), 
        .I2(\vrf/regTable[2][8] ), .I3(\vrf/regTable[3][8] ), .S0(n4929), .S1(
        n4999), .ZN(n3667) );
  MUX4ND0BWP U5485 ( .I0(\vrf/regTable[4][8] ), .I1(\vrf/regTable[5][8] ), 
        .I2(\vrf/regTable[6][8] ), .I3(\vrf/regTable[7][8] ), .S0(n4929), .S1(
        n4999), .ZN(n3668) );
  MUX2D1BWP U5486 ( .I0(n3670), .I1(n3671), .S(n5068), .Z(n3669) );
  MUX4ND0BWP U5487 ( .I0(\vrf/regTable[0][9] ), .I1(\vrf/regTable[1][9] ), 
        .I2(\vrf/regTable[2][9] ), .I3(\vrf/regTable[3][9] ), .S0(n4929), .S1(
        n4999), .ZN(n3670) );
  MUX4ND0BWP U5488 ( .I0(\vrf/regTable[4][9] ), .I1(\vrf/regTable[5][9] ), 
        .I2(\vrf/regTable[6][9] ), .I3(\vrf/regTable[7][9] ), .S0(n4929), .S1(
        n4999), .ZN(n3671) );
  MUX2D1BWP U5489 ( .I0(n3673), .I1(n3674), .S(n5068), .Z(n3672) );
  MUX4ND0BWP U5490 ( .I0(\vrf/regTable[0][10] ), .I1(\vrf/regTable[1][10] ), 
        .I2(\vrf/regTable[2][10] ), .I3(\vrf/regTable[3][10] ), .S0(n4929), 
        .S1(n4999), .ZN(n3673) );
  MUX4ND0BWP U5491 ( .I0(\vrf/regTable[4][10] ), .I1(\vrf/regTable[5][10] ), 
        .I2(\vrf/regTable[6][10] ), .I3(\vrf/regTable[7][10] ), .S0(n4929), 
        .S1(n4999), .ZN(n3674) );
  MUX2D1BWP U5492 ( .I0(n3676), .I1(n3677), .S(n5089), .Z(n3675) );
  MUX4ND0BWP U5493 ( .I0(\srf/regTable[0][0] ), .I1(\srf/regTable[1][0] ), 
        .I2(\srf/regTable[2][0] ), .I3(\srf/regTable[3][0] ), .S0(n4970), .S1(
        n5040), .ZN(n3676) );
  MUX4ND0BWP U5494 ( .I0(\srf/regTable[4][0] ), .I1(\srf/regTable[5][0] ), 
        .I2(\srf/regTable[6][0] ), .I3(\srf/regTable[7][0] ), .S0(n4970), .S1(
        n5040), .ZN(n3677) );
  MUX2D1BWP U5495 ( .I0(n3679), .I1(n3680), .S(n5089), .Z(n3678) );
  MUX4ND0BWP U5496 ( .I0(\srf/regTable[0][1] ), .I1(\srf/regTable[1][1] ), 
        .I2(\srf/regTable[2][1] ), .I3(\srf/regTable[3][1] ), .S0(n4970), .S1(
        n5040), .ZN(n3679) );
  MUX4ND0BWP U5497 ( .I0(\srf/regTable[4][1] ), .I1(\srf/regTable[5][1] ), 
        .I2(\srf/regTable[6][1] ), .I3(\srf/regTable[7][1] ), .S0(n4970), .S1(
        n5040), .ZN(n3680) );
  MUX2D1BWP U5498 ( .I0(n3682), .I1(n3683), .S(n5089), .Z(n3681) );
  MUX4ND0BWP U5499 ( .I0(\srf/regTable[0][2] ), .I1(\srf/regTable[1][2] ), 
        .I2(\srf/regTable[2][2] ), .I3(\srf/regTable[3][2] ), .S0(n4971), .S1(
        n5041), .ZN(n3682) );
  MUX4ND0BWP U5500 ( .I0(\srf/regTable[4][2] ), .I1(\srf/regTable[5][2] ), 
        .I2(\srf/regTable[6][2] ), .I3(\srf/regTable[7][2] ), .S0(n4971), .S1(
        n5041), .ZN(n3683) );
  MUX2D1BWP U5501 ( .I0(n3685), .I1(n3686), .S(n5089), .Z(n3684) );
  MUX4ND0BWP U5502 ( .I0(\srf/regTable[0][5] ), .I1(\srf/regTable[1][5] ), 
        .I2(\srf/regTable[2][5] ), .I3(\srf/regTable[3][5] ), .S0(n4971), .S1(
        n5041), .ZN(n3685) );
  MUX4ND0BWP U5503 ( .I0(\srf/regTable[4][5] ), .I1(\srf/regTable[5][5] ), 
        .I2(\srf/regTable[6][5] ), .I3(\srf/regTable[7][5] ), .S0(n4971), .S1(
        n5041), .ZN(n3686) );
  MUX2D1BWP U5504 ( .I0(n3688), .I1(n3689), .S(n5089), .Z(n3687) );
  MUX4ND0BWP U5505 ( .I0(\srf/regTable[0][6] ), .I1(\srf/regTable[1][6] ), 
        .I2(\srf/regTable[2][6] ), .I3(\srf/regTable[3][6] ), .S0(n4971), .S1(
        n5041), .ZN(n3688) );
  MUX4ND0BWP U5506 ( .I0(\srf/regTable[4][6] ), .I1(\srf/regTable[5][6] ), 
        .I2(\srf/regTable[6][6] ), .I3(\srf/regTable[7][6] ), .S0(n4971), .S1(
        n5041), .ZN(n3689) );
  MUX2D1BWP U5507 ( .I0(n3691), .I1(n3692), .S(n5089), .Z(n3690) );
  MUX4ND0BWP U5508 ( .I0(\srf/regTable[0][7] ), .I1(\srf/regTable[1][7] ), 
        .I2(\srf/regTable[2][7] ), .I3(\srf/regTable[3][7] ), .S0(n4971), .S1(
        n5041), .ZN(n3691) );
  MUX4ND0BWP U5509 ( .I0(\srf/regTable[4][7] ), .I1(\srf/regTable[5][7] ), 
        .I2(\srf/regTable[6][7] ), .I3(\srf/regTable[7][7] ), .S0(n4971), .S1(
        n5041), .ZN(n3692) );
  MUX2D1BWP U5510 ( .I0(n3694), .I1(n3695), .S(n5090), .Z(n3693) );
  MUX4ND0BWP U5511 ( .I0(\srf/regTable[0][8] ), .I1(\srf/regTable[1][8] ), 
        .I2(\srf/regTable[2][8] ), .I3(\srf/regTable[3][8] ), .S0(n4972), .S1(
        n5042), .ZN(n3694) );
  MUX4ND0BWP U5512 ( .I0(\srf/regTable[4][8] ), .I1(\srf/regTable[5][8] ), 
        .I2(\srf/regTable[6][8] ), .I3(\srf/regTable[7][8] ), .S0(n4972), .S1(
        n5042), .ZN(n3695) );
  MUX2D1BWP U5513 ( .I0(n3697), .I1(n3698), .S(n5090), .Z(n3696) );
  MUX4ND0BWP U5514 ( .I0(\srf/regTable[0][9] ), .I1(\srf/regTable[1][9] ), 
        .I2(\srf/regTable[2][9] ), .I3(\srf/regTable[3][9] ), .S0(n4972), .S1(
        n5042), .ZN(n3697) );
  MUX4ND0BWP U5515 ( .I0(\srf/regTable[4][9] ), .I1(\srf/regTable[5][9] ), 
        .I2(\srf/regTable[6][9] ), .I3(\srf/regTable[7][9] ), .S0(n4972), .S1(
        n5042), .ZN(n3698) );
  MUX2D1BWP U5516 ( .I0(n3700), .I1(n3701), .S(n5090), .Z(n3699) );
  MUX4ND0BWP U5517 ( .I0(\srf/regTable[0][10] ), .I1(\srf/regTable[1][10] ), 
        .I2(\srf/regTable[2][10] ), .I3(\srf/regTable[3][10] ), .S0(n4972), 
        .S1(n5042), .ZN(n3700) );
  MUX4ND0BWP U5518 ( .I0(\srf/regTable[4][10] ), .I1(\srf/regTable[5][10] ), 
        .I2(\srf/regTable[6][10] ), .I3(\srf/regTable[7][10] ), .S0(n4972), 
        .S1(n5042), .ZN(n3701) );
  MUX2ND0BWP U5519 ( .I0(n3702), .I1(n3703), .S(n4912), .ZN(vectorData1[239])
         );
  MUX4ND0BWP U5520 ( .I0(\vrf/regTable[0][239] ), .I1(\vrf/regTable[1][239] ), 
        .I2(\vrf/regTable[2][239] ), .I3(\vrf/regTable[3][239] ), .S0(n4792), 
        .S1(n4862), .ZN(n3702) );
  MUX4ND0BWP U5521 ( .I0(\vrf/regTable[4][239] ), .I1(\vrf/regTable[5][239] ), 
        .I2(\vrf/regTable[6][239] ), .I3(\vrf/regTable[7][239] ), .S0(n4792), 
        .S1(n4862), .ZN(n3703) );
  MUX2ND0BWP U5522 ( .I0(n3704), .I1(n3705), .S(n4911), .ZN(vectorData1[224])
         );
  MUX4ND0BWP U5523 ( .I0(\vrf/regTable[0][224] ), .I1(\vrf/regTable[1][224] ), 
        .I2(\vrf/regTable[2][224] ), .I3(\vrf/regTable[3][224] ), .S0(n4790), 
        .S1(n4860), .ZN(n3704) );
  MUX4ND0BWP U5524 ( .I0(\vrf/regTable[4][224] ), .I1(\vrf/regTable[5][224] ), 
        .I2(\vrf/regTable[6][224] ), .I3(\vrf/regTable[7][224] ), .S0(n4790), 
        .S1(n4860), .ZN(n3705) );
  MUX2ND0BWP U5525 ( .I0(n3706), .I1(n3707), .S(n4912), .ZN(vectorData1[238])
         );
  MUX4ND0BWP U5526 ( .I0(\vrf/regTable[0][238] ), .I1(\vrf/regTable[1][238] ), 
        .I2(\vrf/regTable[2][238] ), .I3(\vrf/regTable[3][238] ), .S0(n4792), 
        .S1(n4862), .ZN(n3706) );
  MUX4ND0BWP U5527 ( .I0(\vrf/regTable[4][238] ), .I1(\vrf/regTable[5][238] ), 
        .I2(\vrf/regTable[6][238] ), .I3(\vrf/regTable[7][238] ), .S0(n4792), 
        .S1(n4862), .ZN(n3707) );
  MUX2ND0BWP U5528 ( .I0(n3708), .I1(n3709), .S(n4912), .ZN(vectorData1[237])
         );
  MUX4ND0BWP U5529 ( .I0(\vrf/regTable[0][237] ), .I1(\vrf/regTable[1][237] ), 
        .I2(\vrf/regTable[2][237] ), .I3(\vrf/regTable[3][237] ), .S0(n4792), 
        .S1(n4862), .ZN(n3708) );
  MUX4ND0BWP U5530 ( .I0(\vrf/regTable[4][237] ), .I1(\vrf/regTable[5][237] ), 
        .I2(\vrf/regTable[6][237] ), .I3(\vrf/regTable[7][237] ), .S0(n4792), 
        .S1(n4862), .ZN(n3709) );
  MUX2ND0BWP U5531 ( .I0(n3710), .I1(n3711), .S(n4912), .ZN(vectorData1[236])
         );
  MUX4ND0BWP U5532 ( .I0(\vrf/regTable[0][236] ), .I1(\vrf/regTable[1][236] ), 
        .I2(\vrf/regTable[2][236] ), .I3(\vrf/regTable[3][236] ), .S0(n4792), 
        .S1(n4862), .ZN(n3710) );
  MUX4ND0BWP U5533 ( .I0(\vrf/regTable[4][236] ), .I1(\vrf/regTable[5][236] ), 
        .I2(\vrf/regTable[6][236] ), .I3(\vrf/regTable[7][236] ), .S0(n4792), 
        .S1(n4862), .ZN(n3711) );
  MUX2ND0BWP U5534 ( .I0(n3712), .I1(n3713), .S(n4912), .ZN(vectorData1[235])
         );
  MUX4ND0BWP U5535 ( .I0(\vrf/regTable[0][235] ), .I1(\vrf/regTable[1][235] ), 
        .I2(\vrf/regTable[2][235] ), .I3(\vrf/regTable[3][235] ), .S0(n4792), 
        .S1(n4862), .ZN(n3712) );
  MUX4ND0BWP U5536 ( .I0(\vrf/regTable[4][235] ), .I1(\vrf/regTable[5][235] ), 
        .I2(\vrf/regTable[6][235] ), .I3(\vrf/regTable[7][235] ), .S0(n4792), 
        .S1(n4862), .ZN(n3713) );
  MUX2ND0BWP U5537 ( .I0(n3714), .I1(n3715), .S(n4912), .ZN(vectorData1[234])
         );
  MUX4ND0BWP U5538 ( .I0(\vrf/regTable[0][234] ), .I1(\vrf/regTable[1][234] ), 
        .I2(\vrf/regTable[2][234] ), .I3(\vrf/regTable[3][234] ), .S0(n4792), 
        .S1(n4862), .ZN(n3714) );
  MUX4ND0BWP U5539 ( .I0(\vrf/regTable[4][234] ), .I1(\vrf/regTable[5][234] ), 
        .I2(\vrf/regTable[6][234] ), .I3(\vrf/regTable[7][234] ), .S0(n4792), 
        .S1(n4862), .ZN(n3715) );
  MUX2ND0BWP U5540 ( .I0(n3716), .I1(n3717), .S(n4912), .ZN(vectorData1[233])
         );
  MUX4ND0BWP U5541 ( .I0(\vrf/regTable[0][233] ), .I1(\vrf/regTable[1][233] ), 
        .I2(\vrf/regTable[2][233] ), .I3(\vrf/regTable[3][233] ), .S0(n4791), 
        .S1(n4861), .ZN(n3716) );
  MUX4ND0BWP U5542 ( .I0(\vrf/regTable[4][233] ), .I1(\vrf/regTable[5][233] ), 
        .I2(\vrf/regTable[6][233] ), .I3(\vrf/regTable[7][233] ), .S0(n4791), 
        .S1(n4861), .ZN(n3717) );
  MUX2ND0BWP U5543 ( .I0(n3718), .I1(n3719), .S(n4912), .ZN(vectorData1[232])
         );
  MUX4ND0BWP U5544 ( .I0(\vrf/regTable[0][232] ), .I1(\vrf/regTable[1][232] ), 
        .I2(\vrf/regTable[2][232] ), .I3(\vrf/regTable[3][232] ), .S0(n4791), 
        .S1(n4861), .ZN(n3718) );
  MUX4ND0BWP U5545 ( .I0(\vrf/regTable[4][232] ), .I1(\vrf/regTable[5][232] ), 
        .I2(\vrf/regTable[6][232] ), .I3(\vrf/regTable[7][232] ), .S0(n4791), 
        .S1(n4861), .ZN(n3719) );
  MUX2ND0BWP U5546 ( .I0(n3720), .I1(n3721), .S(n4911), .ZN(vectorData1[225])
         );
  MUX4ND0BWP U5547 ( .I0(\vrf/regTable[0][225] ), .I1(\vrf/regTable[1][225] ), 
        .I2(\vrf/regTable[2][225] ), .I3(\vrf/regTable[3][225] ), .S0(n4790), 
        .S1(n4860), .ZN(n3720) );
  MUX4ND0BWP U5548 ( .I0(\vrf/regTable[4][225] ), .I1(\vrf/regTable[5][225] ), 
        .I2(\vrf/regTable[6][225] ), .I3(\vrf/regTable[7][225] ), .S0(n4790), 
        .S1(n4860), .ZN(n3721) );
  MUX2ND0BWP U5549 ( .I0(n3722), .I1(n3723), .S(n4912), .ZN(vectorData1[231])
         );
  MUX4ND0BWP U5550 ( .I0(\vrf/regTable[0][231] ), .I1(\vrf/regTable[1][231] ), 
        .I2(\vrf/regTable[2][231] ), .I3(\vrf/regTable[3][231] ), .S0(n4791), 
        .S1(n4861), .ZN(n3722) );
  MUX4ND0BWP U5551 ( .I0(\vrf/regTable[4][231] ), .I1(\vrf/regTable[5][231] ), 
        .I2(\vrf/regTable[6][231] ), .I3(\vrf/regTable[7][231] ), .S0(n4791), 
        .S1(n4861), .ZN(n3723) );
  MUX2ND0BWP U5552 ( .I0(n3724), .I1(n3725), .S(n4912), .ZN(vectorData1[230])
         );
  MUX4ND0BWP U5553 ( .I0(\vrf/regTable[0][230] ), .I1(\vrf/regTable[1][230] ), 
        .I2(\vrf/regTable[2][230] ), .I3(\vrf/regTable[3][230] ), .S0(n4791), 
        .S1(n4861), .ZN(n3724) );
  MUX4ND0BWP U5554 ( .I0(\vrf/regTable[4][230] ), .I1(\vrf/regTable[5][230] ), 
        .I2(\vrf/regTable[6][230] ), .I3(\vrf/regTable[7][230] ), .S0(n4791), 
        .S1(n4861), .ZN(n3725) );
  MUX2ND0BWP U5555 ( .I0(n3726), .I1(n3727), .S(n4912), .ZN(vectorData1[229])
         );
  MUX4ND0BWP U5556 ( .I0(\vrf/regTable[0][229] ), .I1(\vrf/regTable[1][229] ), 
        .I2(\vrf/regTable[2][229] ), .I3(\vrf/regTable[3][229] ), .S0(n4791), 
        .S1(n4861), .ZN(n3726) );
  MUX4ND0BWP U5557 ( .I0(\vrf/regTable[4][229] ), .I1(\vrf/regTable[5][229] ), 
        .I2(\vrf/regTable[6][229] ), .I3(\vrf/regTable[7][229] ), .S0(n4791), 
        .S1(n4861), .ZN(n3727) );
  MUX2ND0BWP U5558 ( .I0(n3728), .I1(n3729), .S(n4911), .ZN(vectorData1[226])
         );
  MUX4ND0BWP U5559 ( .I0(\vrf/regTable[0][226] ), .I1(\vrf/regTable[1][226] ), 
        .I2(\vrf/regTable[2][226] ), .I3(\vrf/regTable[3][226] ), .S0(n4790), 
        .S1(n4860), .ZN(n3728) );
  MUX4ND0BWP U5560 ( .I0(\vrf/regTable[4][226] ), .I1(\vrf/regTable[5][226] ), 
        .I2(\vrf/regTable[6][226] ), .I3(\vrf/regTable[7][226] ), .S0(n4790), 
        .S1(n4860), .ZN(n3729) );
  MUX2ND0BWP U5561 ( .I0(n3730), .I1(n3731), .S(n4911), .ZN(vectorData1[227])
         );
  MUX4ND0BWP U5562 ( .I0(\vrf/regTable[0][227] ), .I1(\vrf/regTable[1][227] ), 
        .I2(\vrf/regTable[2][227] ), .I3(\vrf/regTable[3][227] ), .S0(n4790), 
        .S1(n4860), .ZN(n3730) );
  MUX4ND0BWP U5563 ( .I0(\vrf/regTable[4][227] ), .I1(\vrf/regTable[5][227] ), 
        .I2(\vrf/regTable[6][227] ), .I3(\vrf/regTable[7][227] ), .S0(n4790), 
        .S1(n4860), .ZN(n3731) );
  MUX2ND0BWP U5564 ( .I0(n3732), .I1(n3733), .S(n4912), .ZN(vectorData1[228])
         );
  MUX4ND0BWP U5565 ( .I0(\vrf/regTable[0][228] ), .I1(\vrf/regTable[1][228] ), 
        .I2(\vrf/regTable[2][228] ), .I3(\vrf/regTable[3][228] ), .S0(n4791), 
        .S1(n4861), .ZN(n3732) );
  MUX4ND0BWP U5566 ( .I0(\vrf/regTable[4][228] ), .I1(\vrf/regTable[5][228] ), 
        .I2(\vrf/regTable[6][228] ), .I3(\vrf/regTable[7][228] ), .S0(n4791), 
        .S1(n4861), .ZN(n3733) );
  MUX2ND0BWP U5567 ( .I0(n3734), .I1(n3735), .S(n4911), .ZN(vectorData1[223])
         );
  MUX4ND0BWP U5568 ( .I0(\vrf/regTable[0][223] ), .I1(\vrf/regTable[1][223] ), 
        .I2(\vrf/regTable[2][223] ), .I3(\vrf/regTable[3][223] ), .S0(n4790), 
        .S1(n4860), .ZN(n3734) );
  MUX4ND0BWP U5569 ( .I0(\vrf/regTable[4][223] ), .I1(\vrf/regTable[5][223] ), 
        .I2(\vrf/regTable[6][223] ), .I3(\vrf/regTable[7][223] ), .S0(n4790), 
        .S1(n4860), .ZN(n3735) );
  MUX2ND0BWP U5570 ( .I0(n3736), .I1(n3737), .S(n4904), .ZN(vectorData1[143])
         );
  MUX4ND0BWP U5571 ( .I0(\vrf/regTable[0][143] ), .I1(\vrf/regTable[1][143] ), 
        .I2(\vrf/regTable[2][143] ), .I3(\vrf/regTable[3][143] ), .S0(n4776), 
        .S1(n4846), .ZN(n3736) );
  MUX4ND0BWP U5572 ( .I0(\vrf/regTable[4][143] ), .I1(\vrf/regTable[5][143] ), 
        .I2(\vrf/regTable[6][143] ), .I3(\vrf/regTable[7][143] ), .S0(n4776), 
        .S1(n4846), .ZN(n3737) );
  MUX2ND0BWP U5573 ( .I0(n3738), .I1(n3739), .S(n4899), .ZN(vectorData1[79])
         );
  MUX4ND0BWP U5574 ( .I0(\vrf/regTable[0][79] ), .I1(\vrf/regTable[1][79] ), 
        .I2(\vrf/regTable[2][79] ), .I3(\vrf/regTable[3][79] ), .S0(n4766), 
        .S1(n4836), .ZN(n3738) );
  MUX4ND0BWP U5575 ( .I0(\vrf/regTable[4][79] ), .I1(\vrf/regTable[5][79] ), 
        .I2(\vrf/regTable[6][79] ), .I3(\vrf/regTable[7][79] ), .S0(n4766), 
        .S1(n4836), .ZN(n3739) );
  MUX2ND0BWP U5576 ( .I0(n3740), .I1(n3741), .S(n4910), .ZN(vectorData1[207])
         );
  MUX4ND0BWP U5577 ( .I0(\vrf/regTable[0][207] ), .I1(\vrf/regTable[1][207] ), 
        .I2(\vrf/regTable[2][207] ), .I3(\vrf/regTable[3][207] ), .S0(n4787), 
        .S1(n4857), .ZN(n3740) );
  MUX4ND0BWP U5578 ( .I0(\vrf/regTable[4][207] ), .I1(\vrf/regTable[5][207] ), 
        .I2(\vrf/regTable[6][207] ), .I3(\vrf/regTable[7][207] ), .S0(n4787), 
        .S1(n4857), .ZN(n3741) );
  MUX2ND0BWP U5579 ( .I0(n3742), .I1(n3743), .S(n4903), .ZN(vectorData1[128])
         );
  MUX4ND0BWP U5580 ( .I0(\vrf/regTable[0][128] ), .I1(\vrf/regTable[1][128] ), 
        .I2(\vrf/regTable[2][128] ), .I3(\vrf/regTable[3][128] ), .S0(n4774), 
        .S1(n4844), .ZN(n3742) );
  MUX4ND0BWP U5581 ( .I0(\vrf/regTable[4][128] ), .I1(\vrf/regTable[5][128] ), 
        .I2(\vrf/regTable[6][128] ), .I3(\vrf/regTable[7][128] ), .S0(n4774), 
        .S1(n4844), .ZN(n3743) );
  MUX2ND0BWP U5582 ( .I0(n3744), .I1(n3745), .S(n4898), .ZN(vectorData1[64])
         );
  MUX4ND0BWP U5583 ( .I0(\vrf/regTable[0][64] ), .I1(\vrf/regTable[1][64] ), 
        .I2(\vrf/regTable[2][64] ), .I3(\vrf/regTable[3][64] ), .S0(n4763), 
        .S1(n4833), .ZN(n3744) );
  MUX4ND0BWP U5584 ( .I0(\vrf/regTable[4][64] ), .I1(\vrf/regTable[5][64] ), 
        .I2(\vrf/regTable[6][64] ), .I3(\vrf/regTable[7][64] ), .S0(n4763), 
        .S1(n4833), .ZN(n3745) );
  MUX2ND0BWP U5585 ( .I0(n3746), .I1(n3747), .S(n4909), .ZN(vectorData1[192])
         );
  MUX4ND0BWP U5586 ( .I0(\vrf/regTable[0][192] ), .I1(\vrf/regTable[1][192] ), 
        .I2(\vrf/regTable[2][192] ), .I3(\vrf/regTable[3][192] ), .S0(n4785), 
        .S1(n4855), .ZN(n3746) );
  MUX4ND0BWP U5587 ( .I0(\vrf/regTable[4][192] ), .I1(\vrf/regTable[5][192] ), 
        .I2(\vrf/regTable[6][192] ), .I3(\vrf/regTable[7][192] ), .S0(n4785), 
        .S1(n4855), .ZN(n3747) );
  MUX2ND0BWP U5588 ( .I0(n3748), .I1(n3749), .S(n4904), .ZN(vectorData1[142])
         );
  MUX4ND0BWP U5589 ( .I0(\vrf/regTable[0][142] ), .I1(\vrf/regTable[1][142] ), 
        .I2(\vrf/regTable[2][142] ), .I3(\vrf/regTable[3][142] ), .S0(n4776), 
        .S1(n4846), .ZN(n3748) );
  MUX4ND0BWP U5590 ( .I0(\vrf/regTable[4][142] ), .I1(\vrf/regTable[5][142] ), 
        .I2(\vrf/regTable[6][142] ), .I3(\vrf/regTable[7][142] ), .S0(n4776), 
        .S1(n4846), .ZN(n3749) );
  MUX2ND0BWP U5591 ( .I0(n3750), .I1(n3751), .S(n4899), .ZN(vectorData1[78])
         );
  MUX4ND0BWP U5592 ( .I0(\vrf/regTable[0][78] ), .I1(\vrf/regTable[1][78] ), 
        .I2(\vrf/regTable[2][78] ), .I3(\vrf/regTable[3][78] ), .S0(n4766), 
        .S1(n4836), .ZN(n3750) );
  MUX4ND0BWP U5593 ( .I0(\vrf/regTable[4][78] ), .I1(\vrf/regTable[5][78] ), 
        .I2(\vrf/regTable[6][78] ), .I3(\vrf/regTable[7][78] ), .S0(n4766), 
        .S1(n4836), .ZN(n3751) );
  MUX2ND0BWP U5594 ( .I0(n3752), .I1(n3753), .S(n4910), .ZN(vectorData1[206])
         );
  MUX4ND0BWP U5595 ( .I0(\vrf/regTable[0][206] ), .I1(\vrf/regTable[1][206] ), 
        .I2(\vrf/regTable[2][206] ), .I3(\vrf/regTable[3][206] ), .S0(n4787), 
        .S1(n4857), .ZN(n3752) );
  MUX4ND0BWP U5596 ( .I0(\vrf/regTable[4][206] ), .I1(\vrf/regTable[5][206] ), 
        .I2(\vrf/regTable[6][206] ), .I3(\vrf/regTable[7][206] ), .S0(n4787), 
        .S1(n4857), .ZN(n3753) );
  MUX2ND0BWP U5597 ( .I0(n3754), .I1(n3755), .S(n4904), .ZN(vectorData1[141])
         );
  MUX4ND0BWP U5598 ( .I0(\vrf/regTable[0][141] ), .I1(\vrf/regTable[1][141] ), 
        .I2(\vrf/regTable[2][141] ), .I3(\vrf/regTable[3][141] ), .S0(n4776), 
        .S1(n4846), .ZN(n3754) );
  MUX4ND0BWP U5599 ( .I0(\vrf/regTable[4][141] ), .I1(\vrf/regTable[5][141] ), 
        .I2(\vrf/regTable[6][141] ), .I3(\vrf/regTable[7][141] ), .S0(n4776), 
        .S1(n4846), .ZN(n3755) );
  MUX2ND0BWP U5600 ( .I0(n3756), .I1(n3757), .S(n4899), .ZN(vectorData1[77])
         );
  MUX4ND0BWP U5601 ( .I0(\vrf/regTable[0][77] ), .I1(\vrf/regTable[1][77] ), 
        .I2(\vrf/regTable[2][77] ), .I3(\vrf/regTable[3][77] ), .S0(n4765), 
        .S1(n4835), .ZN(n3756) );
  MUX4ND0BWP U5602 ( .I0(\vrf/regTable[4][77] ), .I1(\vrf/regTable[5][77] ), 
        .I2(\vrf/regTable[6][77] ), .I3(\vrf/regTable[7][77] ), .S0(n4765), 
        .S1(n4835), .ZN(n3757) );
  MUX2ND0BWP U5603 ( .I0(n3758), .I1(n3759), .S(n4910), .ZN(vectorData1[205])
         );
  MUX4ND0BWP U5604 ( .I0(\vrf/regTable[0][205] ), .I1(\vrf/regTable[1][205] ), 
        .I2(\vrf/regTable[2][205] ), .I3(\vrf/regTable[3][205] ), .S0(n4787), 
        .S1(n4857), .ZN(n3758) );
  MUX4ND0BWP U5605 ( .I0(\vrf/regTable[4][205] ), .I1(\vrf/regTable[5][205] ), 
        .I2(\vrf/regTable[6][205] ), .I3(\vrf/regTable[7][205] ), .S0(n4787), 
        .S1(n4857), .ZN(n3759) );
  MUX2ND0BWP U5606 ( .I0(n3760), .I1(n3761), .S(n4904), .ZN(vectorData1[140])
         );
  MUX4ND0BWP U5607 ( .I0(\vrf/regTable[0][140] ), .I1(\vrf/regTable[1][140] ), 
        .I2(\vrf/regTable[2][140] ), .I3(\vrf/regTable[3][140] ), .S0(n4776), 
        .S1(n4846), .ZN(n3760) );
  MUX4ND0BWP U5608 ( .I0(\vrf/regTable[4][140] ), .I1(\vrf/regTable[5][140] ), 
        .I2(\vrf/regTable[6][140] ), .I3(\vrf/regTable[7][140] ), .S0(n4776), 
        .S1(n4846), .ZN(n3761) );
  MUX2ND0BWP U5609 ( .I0(n3762), .I1(n3763), .S(n4899), .ZN(vectorData1[76])
         );
  MUX4ND0BWP U5610 ( .I0(\vrf/regTable[0][76] ), .I1(\vrf/regTable[1][76] ), 
        .I2(\vrf/regTable[2][76] ), .I3(\vrf/regTable[3][76] ), .S0(n4765), 
        .S1(n4835), .ZN(n3762) );
  MUX4ND0BWP U5611 ( .I0(\vrf/regTable[4][76] ), .I1(\vrf/regTable[5][76] ), 
        .I2(\vrf/regTable[6][76] ), .I3(\vrf/regTable[7][76] ), .S0(n4765), 
        .S1(n4835), .ZN(n3763) );
  MUX2ND0BWP U5612 ( .I0(n3764), .I1(n3765), .S(n4910), .ZN(vectorData1[204])
         );
  MUX4ND0BWP U5613 ( .I0(\vrf/regTable[0][204] ), .I1(\vrf/regTable[1][204] ), 
        .I2(\vrf/regTable[2][204] ), .I3(\vrf/regTable[3][204] ), .S0(n4787), 
        .S1(n4857), .ZN(n3764) );
  MUX4ND0BWP U5614 ( .I0(\vrf/regTable[4][204] ), .I1(\vrf/regTable[5][204] ), 
        .I2(\vrf/regTable[6][204] ), .I3(\vrf/regTable[7][204] ), .S0(n4787), 
        .S1(n4857), .ZN(n3765) );
  MUX2ND0BWP U5615 ( .I0(n3766), .I1(n3767), .S(n4904), .ZN(vectorData1[139])
         );
  MUX4ND0BWP U5616 ( .I0(\vrf/regTable[0][139] ), .I1(\vrf/regTable[1][139] ), 
        .I2(\vrf/regTable[2][139] ), .I3(\vrf/regTable[3][139] ), .S0(n4776), 
        .S1(n4846), .ZN(n3766) );
  MUX4ND0BWP U5617 ( .I0(\vrf/regTable[4][139] ), .I1(\vrf/regTable[5][139] ), 
        .I2(\vrf/regTable[6][139] ), .I3(\vrf/regTable[7][139] ), .S0(n4776), 
        .S1(n4846), .ZN(n3767) );
  MUX2ND0BWP U5618 ( .I0(n3768), .I1(n3769), .S(n4899), .ZN(vectorData1[75])
         );
  MUX4ND0BWP U5619 ( .I0(\vrf/regTable[0][75] ), .I1(\vrf/regTable[1][75] ), 
        .I2(\vrf/regTable[2][75] ), .I3(\vrf/regTable[3][75] ), .S0(n4765), 
        .S1(n4835), .ZN(n3768) );
  MUX4ND0BWP U5620 ( .I0(\vrf/regTable[4][75] ), .I1(\vrf/regTable[5][75] ), 
        .I2(\vrf/regTable[6][75] ), .I3(\vrf/regTable[7][75] ), .S0(n4765), 
        .S1(n4835), .ZN(n3769) );
  MUX2ND0BWP U5621 ( .I0(n3770), .I1(n3771), .S(n4909), .ZN(vectorData1[203])
         );
  MUX4ND0BWP U5622 ( .I0(\vrf/regTable[0][203] ), .I1(\vrf/regTable[1][203] ), 
        .I2(\vrf/regTable[2][203] ), .I3(\vrf/regTable[3][203] ), .S0(n4786), 
        .S1(n4856), .ZN(n3770) );
  MUX4ND0BWP U5623 ( .I0(\vrf/regTable[4][203] ), .I1(\vrf/regTable[5][203] ), 
        .I2(\vrf/regTable[6][203] ), .I3(\vrf/regTable[7][203] ), .S0(n4786), 
        .S1(n4856), .ZN(n3771) );
  MUX2ND0BWP U5624 ( .I0(n3772), .I1(n3773), .S(n4904), .ZN(vectorData1[138])
         );
  MUX4ND0BWP U5625 ( .I0(\vrf/regTable[0][138] ), .I1(\vrf/regTable[1][138] ), 
        .I2(\vrf/regTable[2][138] ), .I3(\vrf/regTable[3][138] ), .S0(n4776), 
        .S1(n4846), .ZN(n3772) );
  MUX4ND0BWP U5626 ( .I0(\vrf/regTable[4][138] ), .I1(\vrf/regTable[5][138] ), 
        .I2(\vrf/regTable[6][138] ), .I3(\vrf/regTable[7][138] ), .S0(n4776), 
        .S1(n4846), .ZN(n3773) );
  MUX2ND0BWP U5627 ( .I0(n3774), .I1(n3775), .S(n4899), .ZN(vectorData1[74])
         );
  MUX4ND0BWP U5628 ( .I0(\vrf/regTable[0][74] ), .I1(\vrf/regTable[1][74] ), 
        .I2(\vrf/regTable[2][74] ), .I3(\vrf/regTable[3][74] ), .S0(n4765), 
        .S1(n4835), .ZN(n3774) );
  MUX4ND0BWP U5629 ( .I0(\vrf/regTable[4][74] ), .I1(\vrf/regTable[5][74] ), 
        .I2(\vrf/regTable[6][74] ), .I3(\vrf/regTable[7][74] ), .S0(n4765), 
        .S1(n4835), .ZN(n3775) );
  MUX2ND0BWP U5630 ( .I0(n3776), .I1(n3777), .S(n4909), .ZN(vectorData1[202])
         );
  MUX4ND0BWP U5631 ( .I0(\vrf/regTable[0][202] ), .I1(\vrf/regTable[1][202] ), 
        .I2(\vrf/regTable[2][202] ), .I3(\vrf/regTable[3][202] ), .S0(n4786), 
        .S1(n4856), .ZN(n3776) );
  MUX4ND0BWP U5632 ( .I0(\vrf/regTable[4][202] ), .I1(\vrf/regTable[5][202] ), 
        .I2(\vrf/regTable[6][202] ), .I3(\vrf/regTable[7][202] ), .S0(n4786), 
        .S1(n4856), .ZN(n3777) );
  MUX2ND0BWP U5633 ( .I0(n3778), .I1(n3779), .S(n4904), .ZN(vectorData1[137])
         );
  MUX4ND0BWP U5634 ( .I0(\vrf/regTable[0][137] ), .I1(\vrf/regTable[1][137] ), 
        .I2(\vrf/regTable[2][137] ), .I3(\vrf/regTable[3][137] ), .S0(n4775), 
        .S1(n4845), .ZN(n3778) );
  MUX4ND0BWP U5635 ( .I0(\vrf/regTable[4][137] ), .I1(\vrf/regTable[5][137] ), 
        .I2(\vrf/regTable[6][137] ), .I3(\vrf/regTable[7][137] ), .S0(n4775), 
        .S1(n4845), .ZN(n3779) );
  MUX2ND0BWP U5636 ( .I0(n3780), .I1(n3781), .S(n4899), .ZN(vectorData1[73])
         );
  MUX4ND0BWP U5637 ( .I0(\vrf/regTable[0][73] ), .I1(\vrf/regTable[1][73] ), 
        .I2(\vrf/regTable[2][73] ), .I3(\vrf/regTable[3][73] ), .S0(n4765), 
        .S1(n4835), .ZN(n3780) );
  MUX4ND0BWP U5638 ( .I0(\vrf/regTable[4][73] ), .I1(\vrf/regTable[5][73] ), 
        .I2(\vrf/regTable[6][73] ), .I3(\vrf/regTable[7][73] ), .S0(n4765), 
        .S1(n4835), .ZN(n3781) );
  MUX2ND0BWP U5639 ( .I0(n3782), .I1(n3783), .S(n4909), .ZN(vectorData1[201])
         );
  MUX4ND0BWP U5640 ( .I0(\vrf/regTable[0][201] ), .I1(\vrf/regTable[1][201] ), 
        .I2(\vrf/regTable[2][201] ), .I3(\vrf/regTable[3][201] ), .S0(n4786), 
        .S1(n4856), .ZN(n3782) );
  MUX4ND0BWP U5641 ( .I0(\vrf/regTable[4][201] ), .I1(\vrf/regTable[5][201] ), 
        .I2(\vrf/regTable[6][201] ), .I3(\vrf/regTable[7][201] ), .S0(n4786), 
        .S1(n4856), .ZN(n3783) );
  MUX2ND0BWP U5642 ( .I0(n3784), .I1(n3785), .S(n4904), .ZN(vectorData1[136])
         );
  MUX4ND0BWP U5643 ( .I0(\vrf/regTable[0][136] ), .I1(\vrf/regTable[1][136] ), 
        .I2(\vrf/regTable[2][136] ), .I3(\vrf/regTable[3][136] ), .S0(n4775), 
        .S1(n4845), .ZN(n3784) );
  MUX4ND0BWP U5644 ( .I0(\vrf/regTable[4][136] ), .I1(\vrf/regTable[5][136] ), 
        .I2(\vrf/regTable[6][136] ), .I3(\vrf/regTable[7][136] ), .S0(n4775), 
        .S1(n4845), .ZN(n3785) );
  MUX2ND0BWP U5645 ( .I0(n3786), .I1(n3787), .S(n4899), .ZN(vectorData1[72])
         );
  MUX4ND0BWP U5646 ( .I0(\vrf/regTable[0][72] ), .I1(\vrf/regTable[1][72] ), 
        .I2(\vrf/regTable[2][72] ), .I3(\vrf/regTable[3][72] ), .S0(n4765), 
        .S1(n4835), .ZN(n3786) );
  MUX4ND0BWP U5647 ( .I0(\vrf/regTable[4][72] ), .I1(\vrf/regTable[5][72] ), 
        .I2(\vrf/regTable[6][72] ), .I3(\vrf/regTable[7][72] ), .S0(n4765), 
        .S1(n4835), .ZN(n3787) );
  MUX2ND0BWP U5648 ( .I0(n3788), .I1(n3789), .S(n4909), .ZN(vectorData1[200])
         );
  MUX4ND0BWP U5649 ( .I0(\vrf/regTable[0][200] ), .I1(\vrf/regTable[1][200] ), 
        .I2(\vrf/regTable[2][200] ), .I3(\vrf/regTable[3][200] ), .S0(n4786), 
        .S1(n4856), .ZN(n3788) );
  MUX4ND0BWP U5650 ( .I0(\vrf/regTable[4][200] ), .I1(\vrf/regTable[5][200] ), 
        .I2(\vrf/regTable[6][200] ), .I3(\vrf/regTable[7][200] ), .S0(n4786), 
        .S1(n4856), .ZN(n3789) );
  MUX2ND0BWP U5651 ( .I0(n3790), .I1(n3791), .S(n4903), .ZN(vectorData1[129])
         );
  MUX4ND0BWP U5652 ( .I0(\vrf/regTable[0][129] ), .I1(\vrf/regTable[1][129] ), 
        .I2(\vrf/regTable[2][129] ), .I3(\vrf/regTable[3][129] ), .S0(n4774), 
        .S1(n4844), .ZN(n3790) );
  MUX4ND0BWP U5653 ( .I0(\vrf/regTable[4][129] ), .I1(\vrf/regTable[5][129] ), 
        .I2(\vrf/regTable[6][129] ), .I3(\vrf/regTable[7][129] ), .S0(n4774), 
        .S1(n4844), .ZN(n3791) );
  MUX2ND0BWP U5654 ( .I0(n3792), .I1(n3793), .S(n4898), .ZN(vectorData1[65])
         );
  MUX4ND0BWP U5655 ( .I0(\vrf/regTable[0][65] ), .I1(\vrf/regTable[1][65] ), 
        .I2(\vrf/regTable[2][65] ), .I3(\vrf/regTable[3][65] ), .S0(n4763), 
        .S1(n4833), .ZN(n3792) );
  MUX4ND0BWP U5656 ( .I0(\vrf/regTable[4][65] ), .I1(\vrf/regTable[5][65] ), 
        .I2(\vrf/regTable[6][65] ), .I3(\vrf/regTable[7][65] ), .S0(n4763), 
        .S1(n4833), .ZN(n3793) );
  MUX2ND0BWP U5657 ( .I0(n3794), .I1(n3795), .S(n4909), .ZN(vectorData1[193])
         );
  MUX4ND0BWP U5658 ( .I0(\vrf/regTable[0][193] ), .I1(\vrf/regTable[1][193] ), 
        .I2(\vrf/regTable[2][193] ), .I3(\vrf/regTable[3][193] ), .S0(n4785), 
        .S1(n4855), .ZN(n3794) );
  MUX4ND0BWP U5659 ( .I0(\vrf/regTable[4][193] ), .I1(\vrf/regTable[5][193] ), 
        .I2(\vrf/regTable[6][193] ), .I3(\vrf/regTable[7][193] ), .S0(n4785), 
        .S1(n4855), .ZN(n3795) );
  MUX2ND0BWP U5660 ( .I0(n3796), .I1(n3797), .S(n4904), .ZN(vectorData1[135])
         );
  MUX4ND0BWP U5661 ( .I0(\vrf/regTable[0][135] ), .I1(\vrf/regTable[1][135] ), 
        .I2(\vrf/regTable[2][135] ), .I3(\vrf/regTable[3][135] ), .S0(n4775), 
        .S1(n4845), .ZN(n3796) );
  MUX4ND0BWP U5662 ( .I0(\vrf/regTable[4][135] ), .I1(\vrf/regTable[5][135] ), 
        .I2(\vrf/regTable[6][135] ), .I3(\vrf/regTable[7][135] ), .S0(n4775), 
        .S1(n4845), .ZN(n3797) );
  MUX2ND0BWP U5663 ( .I0(n3798), .I1(n3799), .S(n4898), .ZN(vectorData1[71])
         );
  MUX4ND0BWP U5664 ( .I0(\vrf/regTable[0][71] ), .I1(\vrf/regTable[1][71] ), 
        .I2(\vrf/regTable[2][71] ), .I3(\vrf/regTable[3][71] ), .S0(n4764), 
        .S1(n4834), .ZN(n3798) );
  MUX4ND0BWP U5665 ( .I0(\vrf/regTable[4][71] ), .I1(\vrf/regTable[5][71] ), 
        .I2(\vrf/regTable[6][71] ), .I3(\vrf/regTable[7][71] ), .S0(n4764), 
        .S1(n4834), .ZN(n3799) );
  MUX2ND0BWP U5666 ( .I0(n3800), .I1(n3801), .S(n4909), .ZN(vectorData1[199])
         );
  MUX4ND0BWP U5667 ( .I0(\vrf/regTable[0][199] ), .I1(\vrf/regTable[1][199] ), 
        .I2(\vrf/regTable[2][199] ), .I3(\vrf/regTable[3][199] ), .S0(n4786), 
        .S1(n4856), .ZN(n3800) );
  MUX4ND0BWP U5668 ( .I0(\vrf/regTable[4][199] ), .I1(\vrf/regTable[5][199] ), 
        .I2(\vrf/regTable[6][199] ), .I3(\vrf/regTable[7][199] ), .S0(n4786), 
        .S1(n4856), .ZN(n3801) );
  MUX2ND0BWP U5669 ( .I0(n3802), .I1(n3803), .S(n4904), .ZN(vectorData1[134])
         );
  MUX4ND0BWP U5670 ( .I0(\vrf/regTable[0][134] ), .I1(\vrf/regTable[1][134] ), 
        .I2(\vrf/regTable[2][134] ), .I3(\vrf/regTable[3][134] ), .S0(n4775), 
        .S1(n4845), .ZN(n3802) );
  MUX4ND0BWP U5671 ( .I0(\vrf/regTable[4][134] ), .I1(\vrf/regTable[5][134] ), 
        .I2(\vrf/regTable[6][134] ), .I3(\vrf/regTable[7][134] ), .S0(n4775), 
        .S1(n4845), .ZN(n3803) );
  MUX2ND0BWP U5672 ( .I0(n3804), .I1(n3805), .S(n4898), .ZN(vectorData1[70])
         );
  MUX4ND0BWP U5673 ( .I0(\vrf/regTable[0][70] ), .I1(\vrf/regTable[1][70] ), 
        .I2(\vrf/regTable[2][70] ), .I3(\vrf/regTable[3][70] ), .S0(n4764), 
        .S1(n4834), .ZN(n3804) );
  MUX4ND0BWP U5674 ( .I0(\vrf/regTable[4][70] ), .I1(\vrf/regTable[5][70] ), 
        .I2(\vrf/regTable[6][70] ), .I3(\vrf/regTable[7][70] ), .S0(n4764), 
        .S1(n4834), .ZN(n3805) );
  MUX2ND0BWP U5675 ( .I0(n3806), .I1(n3807), .S(n4909), .ZN(vectorData1[198])
         );
  MUX4ND0BWP U5676 ( .I0(\vrf/regTable[0][198] ), .I1(\vrf/regTable[1][198] ), 
        .I2(\vrf/regTable[2][198] ), .I3(\vrf/regTable[3][198] ), .S0(n4786), 
        .S1(n4856), .ZN(n3806) );
  MUX4ND0BWP U5677 ( .I0(\vrf/regTable[4][198] ), .I1(\vrf/regTable[5][198] ), 
        .I2(\vrf/regTable[6][198] ), .I3(\vrf/regTable[7][198] ), .S0(n4786), 
        .S1(n4856), .ZN(n3807) );
  MUX2ND0BWP U5678 ( .I0(n3808), .I1(n3809), .S(n4904), .ZN(vectorData1[133])
         );
  MUX4ND0BWP U5679 ( .I0(\vrf/regTable[0][133] ), .I1(\vrf/regTable[1][133] ), 
        .I2(\vrf/regTable[2][133] ), .I3(\vrf/regTable[3][133] ), .S0(n4775), 
        .S1(n4845), .ZN(n3808) );
  MUX4ND0BWP U5680 ( .I0(\vrf/regTable[4][133] ), .I1(\vrf/regTable[5][133] ), 
        .I2(\vrf/regTable[6][133] ), .I3(\vrf/regTable[7][133] ), .S0(n4775), 
        .S1(n4845), .ZN(n3809) );
  MUX2ND0BWP U5681 ( .I0(n3810), .I1(n3811), .S(n4898), .ZN(vectorData1[69])
         );
  MUX4ND0BWP U5682 ( .I0(\vrf/regTable[0][69] ), .I1(\vrf/regTable[1][69] ), 
        .I2(\vrf/regTable[2][69] ), .I3(\vrf/regTable[3][69] ), .S0(n4764), 
        .S1(n4834), .ZN(n3810) );
  MUX4ND0BWP U5683 ( .I0(\vrf/regTable[4][69] ), .I1(\vrf/regTable[5][69] ), 
        .I2(\vrf/regTable[6][69] ), .I3(\vrf/regTable[7][69] ), .S0(n4764), 
        .S1(n4834), .ZN(n3811) );
  MUX2ND0BWP U5684 ( .I0(n3812), .I1(n3813), .S(n4909), .ZN(vectorData1[197])
         );
  MUX4ND0BWP U5685 ( .I0(\vrf/regTable[0][197] ), .I1(\vrf/regTable[1][197] ), 
        .I2(\vrf/regTable[2][197] ), .I3(\vrf/regTable[3][197] ), .S0(n4785), 
        .S1(n4855), .ZN(n3812) );
  MUX4ND0BWP U5686 ( .I0(\vrf/regTable[4][197] ), .I1(\vrf/regTable[5][197] ), 
        .I2(\vrf/regTable[6][197] ), .I3(\vrf/regTable[7][197] ), .S0(n4785), 
        .S1(n4855), .ZN(n3813) );
  MUX2ND0BWP U5687 ( .I0(n3814), .I1(n3815), .S(n4903), .ZN(vectorData1[130])
         );
  MUX4ND0BWP U5688 ( .I0(\vrf/regTable[0][130] ), .I1(\vrf/regTable[1][130] ), 
        .I2(\vrf/regTable[2][130] ), .I3(\vrf/regTable[3][130] ), .S0(n4774), 
        .S1(n4844), .ZN(n3814) );
  MUX4ND0BWP U5689 ( .I0(\vrf/regTable[4][130] ), .I1(\vrf/regTable[5][130] ), 
        .I2(\vrf/regTable[6][130] ), .I3(\vrf/regTable[7][130] ), .S0(n4774), 
        .S1(n4844), .ZN(n3815) );
  MUX2ND0BWP U5690 ( .I0(n3816), .I1(n3817), .S(n4898), .ZN(vectorData1[66])
         );
  MUX4ND0BWP U5691 ( .I0(\vrf/regTable[0][66] ), .I1(\vrf/regTable[1][66] ), 
        .I2(\vrf/regTable[2][66] ), .I3(\vrf/regTable[3][66] ), .S0(n4764), 
        .S1(n4834), .ZN(n3816) );
  MUX4ND0BWP U5692 ( .I0(\vrf/regTable[4][66] ), .I1(\vrf/regTable[5][66] ), 
        .I2(\vrf/regTable[6][66] ), .I3(\vrf/regTable[7][66] ), .S0(n4764), 
        .S1(n4834), .ZN(n3817) );
  MUX2ND0BWP U5693 ( .I0(n3818), .I1(n3819), .S(n4909), .ZN(vectorData1[194])
         );
  MUX4ND0BWP U5694 ( .I0(\vrf/regTable[0][194] ), .I1(\vrf/regTable[1][194] ), 
        .I2(\vrf/regTable[2][194] ), .I3(\vrf/regTable[3][194] ), .S0(n4785), 
        .S1(n4855), .ZN(n3818) );
  MUX4ND0BWP U5695 ( .I0(\vrf/regTable[4][194] ), .I1(\vrf/regTable[5][194] ), 
        .I2(\vrf/regTable[6][194] ), .I3(\vrf/regTable[7][194] ), .S0(n4785), 
        .S1(n4855), .ZN(n3819) );
  MUX2ND0BWP U5696 ( .I0(n3820), .I1(n3821), .S(n4903), .ZN(vectorData1[131])
         );
  MUX4ND0BWP U5697 ( .I0(\vrf/regTable[0][131] ), .I1(\vrf/regTable[1][131] ), 
        .I2(\vrf/regTable[2][131] ), .I3(\vrf/regTable[3][131] ), .S0(n4774), 
        .S1(n4844), .ZN(n3820) );
  MUX4ND0BWP U5698 ( .I0(\vrf/regTable[4][131] ), .I1(\vrf/regTable[5][131] ), 
        .I2(\vrf/regTable[6][131] ), .I3(\vrf/regTable[7][131] ), .S0(n4774), 
        .S1(n4844), .ZN(n3821) );
  MUX2ND0BWP U5699 ( .I0(n3822), .I1(n3823), .S(n4898), .ZN(vectorData1[67])
         );
  MUX4ND0BWP U5700 ( .I0(\vrf/regTable[0][67] ), .I1(\vrf/regTable[1][67] ), 
        .I2(\vrf/regTable[2][67] ), .I3(\vrf/regTable[3][67] ), .S0(n4764), 
        .S1(n4834), .ZN(n3822) );
  MUX4ND0BWP U5701 ( .I0(\vrf/regTable[4][67] ), .I1(\vrf/regTable[5][67] ), 
        .I2(\vrf/regTable[6][67] ), .I3(\vrf/regTable[7][67] ), .S0(n4764), 
        .S1(n4834), .ZN(n3823) );
  MUX2ND0BWP U5702 ( .I0(n3824), .I1(n3825), .S(n4909), .ZN(vectorData1[195])
         );
  MUX4ND0BWP U5703 ( .I0(\vrf/regTable[0][195] ), .I1(\vrf/regTable[1][195] ), 
        .I2(\vrf/regTable[2][195] ), .I3(\vrf/regTable[3][195] ), .S0(n4785), 
        .S1(n4855), .ZN(n3824) );
  MUX4ND0BWP U5704 ( .I0(\vrf/regTable[4][195] ), .I1(\vrf/regTable[5][195] ), 
        .I2(\vrf/regTable[6][195] ), .I3(\vrf/regTable[7][195] ), .S0(n4785), 
        .S1(n4855), .ZN(n3825) );
  MUX2ND0BWP U5705 ( .I0(n3826), .I1(n3827), .S(n4904), .ZN(vectorData1[132])
         );
  MUX4ND0BWP U5706 ( .I0(\vrf/regTable[0][132] ), .I1(\vrf/regTable[1][132] ), 
        .I2(\vrf/regTable[2][132] ), .I3(\vrf/regTable[3][132] ), .S0(n4775), 
        .S1(n4845), .ZN(n3826) );
  MUX4ND0BWP U5707 ( .I0(\vrf/regTable[4][132] ), .I1(\vrf/regTable[5][132] ), 
        .I2(\vrf/regTable[6][132] ), .I3(\vrf/regTable[7][132] ), .S0(n4775), 
        .S1(n4845), .ZN(n3827) );
  MUX2ND0BWP U5708 ( .I0(n3828), .I1(n3829), .S(n4898), .ZN(vectorData1[68])
         );
  MUX4ND0BWP U5709 ( .I0(\vrf/regTable[0][68] ), .I1(\vrf/regTable[1][68] ), 
        .I2(\vrf/regTable[2][68] ), .I3(\vrf/regTable[3][68] ), .S0(n4764), 
        .S1(n4834), .ZN(n3828) );
  MUX4ND0BWP U5710 ( .I0(\vrf/regTable[4][68] ), .I1(\vrf/regTable[5][68] ), 
        .I2(\vrf/regTable[6][68] ), .I3(\vrf/regTable[7][68] ), .S0(n4764), 
        .S1(n4834), .ZN(n3829) );
  MUX2ND0BWP U5711 ( .I0(n3830), .I1(n3831), .S(n4909), .ZN(vectorData1[196])
         );
  MUX4ND0BWP U5712 ( .I0(\vrf/regTable[0][196] ), .I1(\vrf/regTable[1][196] ), 
        .I2(\vrf/regTable[2][196] ), .I3(\vrf/regTable[3][196] ), .S0(n4785), 
        .S1(n4855), .ZN(n3830) );
  MUX4ND0BWP U5713 ( .I0(\vrf/regTable[4][196] ), .I1(\vrf/regTable[5][196] ), 
        .I2(\vrf/regTable[6][196] ), .I3(\vrf/regTable[7][196] ), .S0(n4785), 
        .S1(n4855), .ZN(n3831) );
  MUX2ND0BWP U5714 ( .I0(n3832), .I1(n3833), .S(n4910), .ZN(vectorData1[208])
         );
  MUX4ND0BWP U5715 ( .I0(\vrf/regTable[0][208] ), .I1(\vrf/regTable[1][208] ), 
        .I2(\vrf/regTable[2][208] ), .I3(\vrf/regTable[3][208] ), .S0(n4787), 
        .S1(n4857), .ZN(n3832) );
  MUX4ND0BWP U5716 ( .I0(\vrf/regTable[4][208] ), .I1(\vrf/regTable[5][208] ), 
        .I2(\vrf/regTable[6][208] ), .I3(\vrf/regTable[7][208] ), .S0(n4787), 
        .S1(n4857), .ZN(n3833) );
  MUX2ND0BWP U5717 ( .I0(n3834), .I1(n3835), .S(n4911), .ZN(vectorData1[222])
         );
  MUX4ND0BWP U5718 ( .I0(\vrf/regTable[0][222] ), .I1(\vrf/regTable[1][222] ), 
        .I2(\vrf/regTable[2][222] ), .I3(\vrf/regTable[3][222] ), .S0(n4790), 
        .S1(n4860), .ZN(n3834) );
  MUX4ND0BWP U5719 ( .I0(\vrf/regTable[4][222] ), .I1(\vrf/regTable[5][222] ), 
        .I2(\vrf/regTable[6][222] ), .I3(\vrf/regTable[7][222] ), .S0(n4790), 
        .S1(n4860), .ZN(n3835) );
  MUX2ND0BWP U5720 ( .I0(n3836), .I1(n3837), .S(n4911), .ZN(vectorData1[221])
         );
  MUX4ND0BWP U5721 ( .I0(\vrf/regTable[0][221] ), .I1(\vrf/regTable[1][221] ), 
        .I2(\vrf/regTable[2][221] ), .I3(\vrf/regTable[3][221] ), .S0(n4789), 
        .S1(n4859), .ZN(n3836) );
  MUX4ND0BWP U5722 ( .I0(\vrf/regTable[4][221] ), .I1(\vrf/regTable[5][221] ), 
        .I2(\vrf/regTable[6][221] ), .I3(\vrf/regTable[7][221] ), .S0(n4789), 
        .S1(n4859), .ZN(n3837) );
  MUX2ND0BWP U5723 ( .I0(n3838), .I1(n3839), .S(n4911), .ZN(vectorData1[220])
         );
  MUX4ND0BWP U5724 ( .I0(\vrf/regTable[0][220] ), .I1(\vrf/regTable[1][220] ), 
        .I2(\vrf/regTable[2][220] ), .I3(\vrf/regTable[3][220] ), .S0(n4789), 
        .S1(n4859), .ZN(n3838) );
  MUX4ND0BWP U5725 ( .I0(\vrf/regTable[4][220] ), .I1(\vrf/regTable[5][220] ), 
        .I2(\vrf/regTable[6][220] ), .I3(\vrf/regTable[7][220] ), .S0(n4789), 
        .S1(n4859), .ZN(n3839) );
  MUX2ND0BWP U5726 ( .I0(n3840), .I1(n3841), .S(n4911), .ZN(vectorData1[219])
         );
  MUX4ND0BWP U5727 ( .I0(\vrf/regTable[0][219] ), .I1(\vrf/regTable[1][219] ), 
        .I2(\vrf/regTable[2][219] ), .I3(\vrf/regTable[3][219] ), .S0(n4789), 
        .S1(n4859), .ZN(n3840) );
  MUX4ND0BWP U5728 ( .I0(\vrf/regTable[4][219] ), .I1(\vrf/regTable[5][219] ), 
        .I2(\vrf/regTable[6][219] ), .I3(\vrf/regTable[7][219] ), .S0(n4789), 
        .S1(n4859), .ZN(n3841) );
  MUX2ND0BWP U5729 ( .I0(n3842), .I1(n3843), .S(n4911), .ZN(vectorData1[218])
         );
  MUX4ND0BWP U5730 ( .I0(\vrf/regTable[0][218] ), .I1(\vrf/regTable[1][218] ), 
        .I2(\vrf/regTable[2][218] ), .I3(\vrf/regTable[3][218] ), .S0(n4789), 
        .S1(n4859), .ZN(n3842) );
  MUX4ND0BWP U5731 ( .I0(\vrf/regTable[4][218] ), .I1(\vrf/regTable[5][218] ), 
        .I2(\vrf/regTable[6][218] ), .I3(\vrf/regTable[7][218] ), .S0(n4789), 
        .S1(n4859), .ZN(n3843) );
  MUX2ND0BWP U5732 ( .I0(n3844), .I1(n3845), .S(n4911), .ZN(vectorData1[217])
         );
  MUX4ND0BWP U5733 ( .I0(\vrf/regTable[0][217] ), .I1(\vrf/regTable[1][217] ), 
        .I2(\vrf/regTable[2][217] ), .I3(\vrf/regTable[3][217] ), .S0(n4789), 
        .S1(n4859), .ZN(n3844) );
  MUX4ND0BWP U5734 ( .I0(\vrf/regTable[4][217] ), .I1(\vrf/regTable[5][217] ), 
        .I2(\vrf/regTable[6][217] ), .I3(\vrf/regTable[7][217] ), .S0(n4789), 
        .S1(n4859), .ZN(n3845) );
  MUX2ND0BWP U5735 ( .I0(n3846), .I1(n3847), .S(n4911), .ZN(vectorData1[216])
         );
  MUX4ND0BWP U5736 ( .I0(\vrf/regTable[0][216] ), .I1(\vrf/regTable[1][216] ), 
        .I2(\vrf/regTable[2][216] ), .I3(\vrf/regTable[3][216] ), .S0(n4789), 
        .S1(n4859), .ZN(n3846) );
  MUX4ND0BWP U5737 ( .I0(\vrf/regTable[4][216] ), .I1(\vrf/regTable[5][216] ), 
        .I2(\vrf/regTable[6][216] ), .I3(\vrf/regTable[7][216] ), .S0(n4789), 
        .S1(n4859), .ZN(n3847) );
  MUX2ND0BWP U5738 ( .I0(n3848), .I1(n3849), .S(n4910), .ZN(vectorData1[209])
         );
  MUX4ND0BWP U5739 ( .I0(\vrf/regTable[0][209] ), .I1(\vrf/regTable[1][209] ), 
        .I2(\vrf/regTable[2][209] ), .I3(\vrf/regTable[3][209] ), .S0(n4787), 
        .S1(n4857), .ZN(n3848) );
  MUX4ND0BWP U5740 ( .I0(\vrf/regTable[4][209] ), .I1(\vrf/regTable[5][209] ), 
        .I2(\vrf/regTable[6][209] ), .I3(\vrf/regTable[7][209] ), .S0(n4787), 
        .S1(n4857), .ZN(n3849) );
  MUX2ND0BWP U5741 ( .I0(n3850), .I1(n3851), .S(n4910), .ZN(vectorData1[215])
         );
  MUX4ND0BWP U5742 ( .I0(\vrf/regTable[0][215] ), .I1(\vrf/regTable[1][215] ), 
        .I2(\vrf/regTable[2][215] ), .I3(\vrf/regTable[3][215] ), .S0(n4788), 
        .S1(n4858), .ZN(n3850) );
  MUX4ND0BWP U5743 ( .I0(\vrf/regTable[4][215] ), .I1(\vrf/regTable[5][215] ), 
        .I2(\vrf/regTable[6][215] ), .I3(\vrf/regTable[7][215] ), .S0(n4788), 
        .S1(n4858), .ZN(n3851) );
  MUX2ND0BWP U5744 ( .I0(n3852), .I1(n3853), .S(n4910), .ZN(vectorData1[214])
         );
  MUX4ND0BWP U5745 ( .I0(\vrf/regTable[0][214] ), .I1(\vrf/regTable[1][214] ), 
        .I2(\vrf/regTable[2][214] ), .I3(\vrf/regTable[3][214] ), .S0(n4788), 
        .S1(n4858), .ZN(n3852) );
  MUX4ND0BWP U5746 ( .I0(\vrf/regTable[4][214] ), .I1(\vrf/regTable[5][214] ), 
        .I2(\vrf/regTable[6][214] ), .I3(\vrf/regTable[7][214] ), .S0(n4788), 
        .S1(n4858), .ZN(n3853) );
  MUX2ND0BWP U5747 ( .I0(n3854), .I1(n3855), .S(n4910), .ZN(vectorData1[213])
         );
  MUX4ND0BWP U5748 ( .I0(\vrf/regTable[0][213] ), .I1(\vrf/regTable[1][213] ), 
        .I2(\vrf/regTable[2][213] ), .I3(\vrf/regTable[3][213] ), .S0(n4788), 
        .S1(n4858), .ZN(n3854) );
  MUX4ND0BWP U5749 ( .I0(\vrf/regTable[4][213] ), .I1(\vrf/regTable[5][213] ), 
        .I2(\vrf/regTable[6][213] ), .I3(\vrf/regTable[7][213] ), .S0(n4788), 
        .S1(n4858), .ZN(n3855) );
  MUX2ND0BWP U5750 ( .I0(n3856), .I1(n3857), .S(n4910), .ZN(vectorData1[210])
         );
  MUX4ND0BWP U5751 ( .I0(\vrf/regTable[0][210] ), .I1(\vrf/regTable[1][210] ), 
        .I2(\vrf/regTable[2][210] ), .I3(\vrf/regTable[3][210] ), .S0(n4788), 
        .S1(n4858), .ZN(n3856) );
  MUX4ND0BWP U5752 ( .I0(\vrf/regTable[4][210] ), .I1(\vrf/regTable[5][210] ), 
        .I2(\vrf/regTable[6][210] ), .I3(\vrf/regTable[7][210] ), .S0(n4788), 
        .S1(n4858), .ZN(n3857) );
  MUX2ND0BWP U5753 ( .I0(n3858), .I1(n3859), .S(n4910), .ZN(vectorData1[211])
         );
  MUX4ND0BWP U5754 ( .I0(\vrf/regTable[0][211] ), .I1(\vrf/regTable[1][211] ), 
        .I2(\vrf/regTable[2][211] ), .I3(\vrf/regTable[3][211] ), .S0(n4788), 
        .S1(n4858), .ZN(n3858) );
  MUX4ND0BWP U5755 ( .I0(\vrf/regTable[4][211] ), .I1(\vrf/regTable[5][211] ), 
        .I2(\vrf/regTable[6][211] ), .I3(\vrf/regTable[7][211] ), .S0(n4788), 
        .S1(n4858), .ZN(n3859) );
  MUX2ND0BWP U5756 ( .I0(n3860), .I1(n3861), .S(n4910), .ZN(vectorData1[212])
         );
  MUX4ND0BWP U5757 ( .I0(\vrf/regTable[0][212] ), .I1(\vrf/regTable[1][212] ), 
        .I2(\vrf/regTable[2][212] ), .I3(\vrf/regTable[3][212] ), .S0(n4788), 
        .S1(n4858), .ZN(n3860) );
  MUX4ND0BWP U5758 ( .I0(\vrf/regTable[4][212] ), .I1(\vrf/regTable[5][212] ), 
        .I2(\vrf/regTable[6][212] ), .I3(\vrf/regTable[7][212] ), .S0(n4788), 
        .S1(n4858), .ZN(n3861) );
  MUX2ND0BWP U5759 ( .I0(n3862), .I1(n3863), .S(n4914), .ZN(vectorData1[255])
         );
  MUX4ND0BWP U5760 ( .I0(\vrf/regTable[0][255] ), .I1(\vrf/regTable[1][255] ), 
        .I2(\vrf/regTable[2][255] ), .I3(\vrf/regTable[3][255] ), .S0(n4795), 
        .S1(n4865), .ZN(n3862) );
  MUX4ND0BWP U5761 ( .I0(\vrf/regTable[4][255] ), .I1(\vrf/regTable[5][255] ), 
        .I2(\vrf/regTable[6][255] ), .I3(\vrf/regTable[7][255] ), .S0(n4795), 
        .S1(n4865), .ZN(n3863) );
  MUX2ND0BWP U5762 ( .I0(n3864), .I1(n3865), .S(n4913), .ZN(vectorData1[240])
         );
  MUX4ND0BWP U5763 ( .I0(\vrf/regTable[0][240] ), .I1(\vrf/regTable[1][240] ), 
        .I2(\vrf/regTable[2][240] ), .I3(\vrf/regTable[3][240] ), .S0(n4793), 
        .S1(n4863), .ZN(n3864) );
  MUX4ND0BWP U5764 ( .I0(\vrf/regTable[4][240] ), .I1(\vrf/regTable[5][240] ), 
        .I2(\vrf/regTable[6][240] ), .I3(\vrf/regTable[7][240] ), .S0(n4793), 
        .S1(n4863), .ZN(n3865) );
  MUX2ND0BWP U5765 ( .I0(n3866), .I1(n3867), .S(n4914), .ZN(vectorData1[254])
         );
  MUX4ND0BWP U5766 ( .I0(\vrf/regTable[0][254] ), .I1(\vrf/regTable[1][254] ), 
        .I2(\vrf/regTable[2][254] ), .I3(\vrf/regTable[3][254] ), .S0(n4795), 
        .S1(n4865), .ZN(n3866) );
  MUX4ND0BWP U5767 ( .I0(\vrf/regTable[4][254] ), .I1(\vrf/regTable[5][254] ), 
        .I2(\vrf/regTable[6][254] ), .I3(\vrf/regTable[7][254] ), .S0(n4795), 
        .S1(n4865), .ZN(n3867) );
  MUX2ND0BWP U5768 ( .I0(n3868), .I1(n3869), .S(n4914), .ZN(vectorData1[253])
         );
  MUX4ND0BWP U5769 ( .I0(\vrf/regTable[0][253] ), .I1(\vrf/regTable[1][253] ), 
        .I2(\vrf/regTable[2][253] ), .I3(\vrf/regTable[3][253] ), .S0(n4795), 
        .S1(n4865), .ZN(n3868) );
  MUX4ND0BWP U5770 ( .I0(\vrf/regTable[4][253] ), .I1(\vrf/regTable[5][253] ), 
        .I2(\vrf/regTable[6][253] ), .I3(\vrf/regTable[7][253] ), .S0(n4795), 
        .S1(n4865), .ZN(n3869) );
  MUX2ND0BWP U5771 ( .I0(n3870), .I1(n3871), .S(n4914), .ZN(vectorData1[252])
         );
  MUX4ND0BWP U5772 ( .I0(\vrf/regTable[0][252] ), .I1(\vrf/regTable[1][252] ), 
        .I2(\vrf/regTable[2][252] ), .I3(\vrf/regTable[3][252] ), .S0(n4795), 
        .S1(n4865), .ZN(n3870) );
  MUX4ND0BWP U5773 ( .I0(\vrf/regTable[4][252] ), .I1(\vrf/regTable[5][252] ), 
        .I2(\vrf/regTable[6][252] ), .I3(\vrf/regTable[7][252] ), .S0(n4795), 
        .S1(n4865), .ZN(n3871) );
  MUX2ND0BWP U5774 ( .I0(n3872), .I1(n3873), .S(n4913), .ZN(vectorData1[251])
         );
  MUX4ND0BWP U5775 ( .I0(\vrf/regTable[0][251] ), .I1(\vrf/regTable[1][251] ), 
        .I2(\vrf/regTable[2][251] ), .I3(\vrf/regTable[3][251] ), .S0(n4794), 
        .S1(n4864), .ZN(n3872) );
  MUX4ND0BWP U5776 ( .I0(\vrf/regTable[4][251] ), .I1(\vrf/regTable[5][251] ), 
        .I2(\vrf/regTable[6][251] ), .I3(\vrf/regTable[7][251] ), .S0(n4794), 
        .S1(n4864), .ZN(n3873) );
  MUX2ND0BWP U5777 ( .I0(n3874), .I1(n3875), .S(n4913), .ZN(vectorData1[250])
         );
  MUX4ND0BWP U5778 ( .I0(\vrf/regTable[0][250] ), .I1(\vrf/regTable[1][250] ), 
        .I2(\vrf/regTable[2][250] ), .I3(\vrf/regTable[3][250] ), .S0(n4794), 
        .S1(n4864), .ZN(n3874) );
  MUX4ND0BWP U5779 ( .I0(\vrf/regTable[4][250] ), .I1(\vrf/regTable[5][250] ), 
        .I2(\vrf/regTable[6][250] ), .I3(\vrf/regTable[7][250] ), .S0(n4794), 
        .S1(n4864), .ZN(n3875) );
  MUX2ND0BWP U5780 ( .I0(n3876), .I1(n3877), .S(n4913), .ZN(vectorData1[249])
         );
  MUX4ND0BWP U5781 ( .I0(\vrf/regTable[0][249] ), .I1(\vrf/regTable[1][249] ), 
        .I2(\vrf/regTable[2][249] ), .I3(\vrf/regTable[3][249] ), .S0(n4794), 
        .S1(n4864), .ZN(n3876) );
  MUX4ND0BWP U5782 ( .I0(\vrf/regTable[4][249] ), .I1(\vrf/regTable[5][249] ), 
        .I2(\vrf/regTable[6][249] ), .I3(\vrf/regTable[7][249] ), .S0(n4794), 
        .S1(n4864), .ZN(n3877) );
  MUX2ND0BWP U5783 ( .I0(n3878), .I1(n3879), .S(n4913), .ZN(vectorData1[248])
         );
  MUX4ND0BWP U5784 ( .I0(\vrf/regTable[0][248] ), .I1(\vrf/regTable[1][248] ), 
        .I2(\vrf/regTable[2][248] ), .I3(\vrf/regTable[3][248] ), .S0(n4794), 
        .S1(n4864), .ZN(n3878) );
  MUX4ND0BWP U5785 ( .I0(\vrf/regTable[4][248] ), .I1(\vrf/regTable[5][248] ), 
        .I2(\vrf/regTable[6][248] ), .I3(\vrf/regTable[7][248] ), .S0(n4794), 
        .S1(n4864), .ZN(n3879) );
  MUX2ND0BWP U5786 ( .I0(n3880), .I1(n3881), .S(n4913), .ZN(vectorData1[241])
         );
  MUX4ND0BWP U5787 ( .I0(\vrf/regTable[0][241] ), .I1(\vrf/regTable[1][241] ), 
        .I2(\vrf/regTable[2][241] ), .I3(\vrf/regTable[3][241] ), .S0(n4793), 
        .S1(n4863), .ZN(n3880) );
  MUX4ND0BWP U5788 ( .I0(\vrf/regTable[4][241] ), .I1(\vrf/regTable[5][241] ), 
        .I2(\vrf/regTable[6][241] ), .I3(\vrf/regTable[7][241] ), .S0(n4793), 
        .S1(n4863), .ZN(n3881) );
  MUX2ND0BWP U5789 ( .I0(n3882), .I1(n3883), .S(n4913), .ZN(vectorData1[247])
         );
  MUX4ND0BWP U5790 ( .I0(\vrf/regTable[0][247] ), .I1(\vrf/regTable[1][247] ), 
        .I2(\vrf/regTable[2][247] ), .I3(\vrf/regTable[3][247] ), .S0(n4794), 
        .S1(n4864), .ZN(n3882) );
  MUX4ND0BWP U5791 ( .I0(\vrf/regTable[4][247] ), .I1(\vrf/regTable[5][247] ), 
        .I2(\vrf/regTable[6][247] ), .I3(\vrf/regTable[7][247] ), .S0(n4794), 
        .S1(n4864), .ZN(n3883) );
  MUX2ND0BWP U5792 ( .I0(n3884), .I1(n3885), .S(n4913), .ZN(vectorData1[246])
         );
  MUX4ND0BWP U5793 ( .I0(\vrf/regTable[0][246] ), .I1(\vrf/regTable[1][246] ), 
        .I2(\vrf/regTable[2][246] ), .I3(\vrf/regTable[3][246] ), .S0(n4794), 
        .S1(n4864), .ZN(n3884) );
  MUX4ND0BWP U5794 ( .I0(\vrf/regTable[4][246] ), .I1(\vrf/regTable[5][246] ), 
        .I2(\vrf/regTable[6][246] ), .I3(\vrf/regTable[7][246] ), .S0(n4794), 
        .S1(n4864), .ZN(n3885) );
  MUX2ND0BWP U5795 ( .I0(n3886), .I1(n3887), .S(n4913), .ZN(vectorData1[245])
         );
  MUX4ND0BWP U5796 ( .I0(\vrf/regTable[0][245] ), .I1(\vrf/regTable[1][245] ), 
        .I2(\vrf/regTable[2][245] ), .I3(\vrf/regTable[3][245] ), .S0(n4793), 
        .S1(n4863), .ZN(n3886) );
  MUX4ND0BWP U5797 ( .I0(\vrf/regTable[4][245] ), .I1(\vrf/regTable[5][245] ), 
        .I2(\vrf/regTable[6][245] ), .I3(\vrf/regTable[7][245] ), .S0(n4793), 
        .S1(n4863), .ZN(n3887) );
  MUX2ND0BWP U5798 ( .I0(n3888), .I1(n3889), .S(n4913), .ZN(vectorData1[242])
         );
  MUX4ND0BWP U5799 ( .I0(\vrf/regTable[0][242] ), .I1(\vrf/regTable[1][242] ), 
        .I2(\vrf/regTable[2][242] ), .I3(\vrf/regTable[3][242] ), .S0(n4793), 
        .S1(n4863), .ZN(n3888) );
  MUX4ND0BWP U5800 ( .I0(\vrf/regTable[4][242] ), .I1(\vrf/regTable[5][242] ), 
        .I2(\vrf/regTable[6][242] ), .I3(\vrf/regTable[7][242] ), .S0(n4793), 
        .S1(n4863), .ZN(n3889) );
  MUX2ND0BWP U5801 ( .I0(n3890), .I1(n3891), .S(n4913), .ZN(vectorData1[243])
         );
  MUX4ND0BWP U5802 ( .I0(\vrf/regTable[0][243] ), .I1(\vrf/regTable[1][243] ), 
        .I2(\vrf/regTable[2][243] ), .I3(\vrf/regTable[3][243] ), .S0(n4793), 
        .S1(n4863), .ZN(n3890) );
  MUX4ND0BWP U5803 ( .I0(\vrf/regTable[4][243] ), .I1(\vrf/regTable[5][243] ), 
        .I2(\vrf/regTable[6][243] ), .I3(\vrf/regTable[7][243] ), .S0(n4793), 
        .S1(n4863), .ZN(n3891) );
  MUX2ND0BWP U5804 ( .I0(n3892), .I1(n3893), .S(n4913), .ZN(vectorData1[244])
         );
  MUX4ND0BWP U5805 ( .I0(\vrf/regTable[0][244] ), .I1(\vrf/regTable[1][244] ), 
        .I2(\vrf/regTable[2][244] ), .I3(\vrf/regTable[3][244] ), .S0(n4793), 
        .S1(n4863), .ZN(n3892) );
  MUX4ND0BWP U5806 ( .I0(\vrf/regTable[4][244] ), .I1(\vrf/regTable[5][244] ), 
        .I2(\vrf/regTable[6][244] ), .I3(\vrf/regTable[7][244] ), .S0(n4793), 
        .S1(n4863), .ZN(n3893) );
  MUX2ND0BWP U5807 ( .I0(n3894), .I1(n3895), .S(n4903), .ZN(vectorData1[127])
         );
  MUX4ND0BWP U5808 ( .I0(\vrf/regTable[0][127] ), .I1(\vrf/regTable[1][127] ), 
        .I2(\vrf/regTable[2][127] ), .I3(\vrf/regTable[3][127] ), .S0(n4774), 
        .S1(n4844), .ZN(n3894) );
  MUX4ND0BWP U5809 ( .I0(\vrf/regTable[4][127] ), .I1(\vrf/regTable[5][127] ), 
        .I2(\vrf/regTable[6][127] ), .I3(\vrf/regTable[7][127] ), .S0(n4774), 
        .S1(n4844), .ZN(n3895) );
  MUX2ND0BWP U5810 ( .I0(n3896), .I1(n3897), .S(n4898), .ZN(vectorData1[63])
         );
  MUX4ND0BWP U5811 ( .I0(\vrf/regTable[0][63] ), .I1(\vrf/regTable[1][63] ), 
        .I2(\vrf/regTable[2][63] ), .I3(\vrf/regTable[3][63] ), .S0(n4763), 
        .S1(n4833), .ZN(n3896) );
  MUX4ND0BWP U5812 ( .I0(\vrf/regTable[4][63] ), .I1(\vrf/regTable[5][63] ), 
        .I2(\vrf/regTable[6][63] ), .I3(\vrf/regTable[7][63] ), .S0(n4763), 
        .S1(n4833), .ZN(n3897) );
  MUX2ND0BWP U5813 ( .I0(n3898), .I1(n3899), .S(n4908), .ZN(vectorData1[191])
         );
  MUX4ND0BWP U5814 ( .I0(\vrf/regTable[0][191] ), .I1(\vrf/regTable[1][191] ), 
        .I2(\vrf/regTable[2][191] ), .I3(\vrf/regTable[3][191] ), .S0(n4784), 
        .S1(n4854), .ZN(n3898) );
  MUX4ND0BWP U5815 ( .I0(\vrf/regTable[4][191] ), .I1(\vrf/regTable[5][191] ), 
        .I2(\vrf/regTable[6][191] ), .I3(\vrf/regTable[7][191] ), .S0(n4784), 
        .S1(n4854), .ZN(n3899) );
  MUX2ND0BWP U5816 ( .I0(n3900), .I1(n3901), .S(n4902), .ZN(vectorData1[112])
         );
  MUX4ND0BWP U5817 ( .I0(\vrf/regTable[0][112] ), .I1(\vrf/regTable[1][112] ), 
        .I2(\vrf/regTable[2][112] ), .I3(\vrf/regTable[3][112] ), .S0(n4771), 
        .S1(n4841), .ZN(n3900) );
  MUX4ND0BWP U5818 ( .I0(\vrf/regTable[4][112] ), .I1(\vrf/regTable[5][112] ), 
        .I2(\vrf/regTable[6][112] ), .I3(\vrf/regTable[7][112] ), .S0(n4771), 
        .S1(n4841), .ZN(n3901) );
  MUX2ND0BWP U5819 ( .I0(n3902), .I1(n3903), .S(n4897), .ZN(vectorData1[48])
         );
  MUX4ND0BWP U5820 ( .I0(\vrf/regTable[0][48] ), .I1(\vrf/regTable[1][48] ), 
        .I2(\vrf/regTable[2][48] ), .I3(\vrf/regTable[3][48] ), .S0(n4761), 
        .S1(n4831), .ZN(n3902) );
  MUX4ND0BWP U5821 ( .I0(\vrf/regTable[4][48] ), .I1(\vrf/regTable[5][48] ), 
        .I2(\vrf/regTable[6][48] ), .I3(\vrf/regTable[7][48] ), .S0(n4761), 
        .S1(n4831), .ZN(n3903) );
  MUX2ND0BWP U5822 ( .I0(n3904), .I1(n3905), .S(n4907), .ZN(vectorData1[176])
         );
  MUX4ND0BWP U5823 ( .I0(\vrf/regTable[0][176] ), .I1(\vrf/regTable[1][176] ), 
        .I2(\vrf/regTable[2][176] ), .I3(\vrf/regTable[3][176] ), .S0(n4782), 
        .S1(n4852), .ZN(n3904) );
  MUX4ND0BWP U5824 ( .I0(\vrf/regTable[4][176] ), .I1(\vrf/regTable[5][176] ), 
        .I2(\vrf/regTable[6][176] ), .I3(\vrf/regTable[7][176] ), .S0(n4782), 
        .S1(n4852), .ZN(n3905) );
  MUX2ND0BWP U5825 ( .I0(n3906), .I1(n3907), .S(n4903), .ZN(vectorData1[126])
         );
  MUX4ND0BWP U5826 ( .I0(\vrf/regTable[0][126] ), .I1(\vrf/regTable[1][126] ), 
        .I2(\vrf/regTable[2][126] ), .I3(\vrf/regTable[3][126] ), .S0(n4774), 
        .S1(n4844), .ZN(n3906) );
  MUX4ND0BWP U5827 ( .I0(\vrf/regTable[4][126] ), .I1(\vrf/regTable[5][126] ), 
        .I2(\vrf/regTable[6][126] ), .I3(\vrf/regTable[7][126] ), .S0(n4774), 
        .S1(n4844), .ZN(n3907) );
  MUX2ND0BWP U5828 ( .I0(n3908), .I1(n3909), .S(n4898), .ZN(vectorData1[62])
         );
  MUX4ND0BWP U5829 ( .I0(\vrf/regTable[0][62] ), .I1(\vrf/regTable[1][62] ), 
        .I2(\vrf/regTable[2][62] ), .I3(\vrf/regTable[3][62] ), .S0(n4763), 
        .S1(n4833), .ZN(n3908) );
  MUX4ND0BWP U5830 ( .I0(\vrf/regTable[4][62] ), .I1(\vrf/regTable[5][62] ), 
        .I2(\vrf/regTable[6][62] ), .I3(\vrf/regTable[7][62] ), .S0(n4763), 
        .S1(n4833), .ZN(n3909) );
  MUX2ND0BWP U5831 ( .I0(n3910), .I1(n3911), .S(n4908), .ZN(vectorData1[190])
         );
  MUX4ND0BWP U5832 ( .I0(\vrf/regTable[0][190] ), .I1(\vrf/regTable[1][190] ), 
        .I2(\vrf/regTable[2][190] ), .I3(\vrf/regTable[3][190] ), .S0(n4784), 
        .S1(n4854), .ZN(n3910) );
  MUX4ND0BWP U5833 ( .I0(\vrf/regTable[4][190] ), .I1(\vrf/regTable[5][190] ), 
        .I2(\vrf/regTable[6][190] ), .I3(\vrf/regTable[7][190] ), .S0(n4784), 
        .S1(n4854), .ZN(n3911) );
  MUX2ND0BWP U5834 ( .I0(n3912), .I1(n3913), .S(n4903), .ZN(vectorData1[125])
         );
  MUX4ND0BWP U5835 ( .I0(\vrf/regTable[0][125] ), .I1(\vrf/regTable[1][125] ), 
        .I2(\vrf/regTable[2][125] ), .I3(\vrf/regTable[3][125] ), .S0(n4773), 
        .S1(n4843), .ZN(n3912) );
  MUX4ND0BWP U5836 ( .I0(\vrf/regTable[4][125] ), .I1(\vrf/regTable[5][125] ), 
        .I2(\vrf/regTable[6][125] ), .I3(\vrf/regTable[7][125] ), .S0(n4773), 
        .S1(n4843), .ZN(n3913) );
  MUX2ND0BWP U5837 ( .I0(n3914), .I1(n3915), .S(n4898), .ZN(vectorData1[61])
         );
  MUX4ND0BWP U5838 ( .I0(\vrf/regTable[0][61] ), .I1(\vrf/regTable[1][61] ), 
        .I2(\vrf/regTable[2][61] ), .I3(\vrf/regTable[3][61] ), .S0(n4763), 
        .S1(n4833), .ZN(n3914) );
  MUX4ND0BWP U5839 ( .I0(\vrf/regTable[4][61] ), .I1(\vrf/regTable[5][61] ), 
        .I2(\vrf/regTable[6][61] ), .I3(\vrf/regTable[7][61] ), .S0(n4763), 
        .S1(n4833), .ZN(n3915) );
  MUX2ND0BWP U5840 ( .I0(n3916), .I1(n3917), .S(n4908), .ZN(vectorData1[189])
         );
  MUX4ND0BWP U5841 ( .I0(\vrf/regTable[0][189] ), .I1(\vrf/regTable[1][189] ), 
        .I2(\vrf/regTable[2][189] ), .I3(\vrf/regTable[3][189] ), .S0(n4784), 
        .S1(n4854), .ZN(n3916) );
  MUX4ND0BWP U5842 ( .I0(\vrf/regTable[4][189] ), .I1(\vrf/regTable[5][189] ), 
        .I2(\vrf/regTable[6][189] ), .I3(\vrf/regTable[7][189] ), .S0(n4784), 
        .S1(n4854), .ZN(n3917) );
  MUX2ND0BWP U5843 ( .I0(n3918), .I1(n3919), .S(n4903), .ZN(vectorData1[124])
         );
  MUX4ND0BWP U5844 ( .I0(\vrf/regTable[0][124] ), .I1(\vrf/regTable[1][124] ), 
        .I2(\vrf/regTable[2][124] ), .I3(\vrf/regTable[3][124] ), .S0(n4773), 
        .S1(n4843), .ZN(n3918) );
  MUX4ND0BWP U5845 ( .I0(\vrf/regTable[4][124] ), .I1(\vrf/regTable[5][124] ), 
        .I2(\vrf/regTable[6][124] ), .I3(\vrf/regTable[7][124] ), .S0(n4773), 
        .S1(n4843), .ZN(n3919) );
  MUX2ND0BWP U5846 ( .I0(n3920), .I1(n3921), .S(n4898), .ZN(vectorData1[60])
         );
  MUX4ND0BWP U5847 ( .I0(\vrf/regTable[0][60] ), .I1(\vrf/regTable[1][60] ), 
        .I2(\vrf/regTable[2][60] ), .I3(\vrf/regTable[3][60] ), .S0(n4763), 
        .S1(n4833), .ZN(n3920) );
  MUX4ND0BWP U5848 ( .I0(\vrf/regTable[4][60] ), .I1(\vrf/regTable[5][60] ), 
        .I2(\vrf/regTable[6][60] ), .I3(\vrf/regTable[7][60] ), .S0(n4763), 
        .S1(n4833), .ZN(n3921) );
  MUX2ND0BWP U5849 ( .I0(n3922), .I1(n3923), .S(n4908), .ZN(vectorData1[188])
         );
  MUX4ND0BWP U5850 ( .I0(\vrf/regTable[0][188] ), .I1(\vrf/regTable[1][188] ), 
        .I2(\vrf/regTable[2][188] ), .I3(\vrf/regTable[3][188] ), .S0(n4784), 
        .S1(n4854), .ZN(n3922) );
  MUX4ND0BWP U5851 ( .I0(\vrf/regTable[4][188] ), .I1(\vrf/regTable[5][188] ), 
        .I2(\vrf/regTable[6][188] ), .I3(\vrf/regTable[7][188] ), .S0(n4784), 
        .S1(n4854), .ZN(n3923) );
  MUX2ND0BWP U5852 ( .I0(n3924), .I1(n3925), .S(n4903), .ZN(vectorData1[123])
         );
  MUX4ND0BWP U5853 ( .I0(\vrf/regTable[0][123] ), .I1(\vrf/regTable[1][123] ), 
        .I2(\vrf/regTable[2][123] ), .I3(\vrf/regTable[3][123] ), .S0(n4773), 
        .S1(n4843), .ZN(n3924) );
  MUX4ND0BWP U5854 ( .I0(\vrf/regTable[4][123] ), .I1(\vrf/regTable[5][123] ), 
        .I2(\vrf/regTable[6][123] ), .I3(\vrf/regTable[7][123] ), .S0(n4773), 
        .S1(n4843), .ZN(n3925) );
  MUX2ND0BWP U5855 ( .I0(n3926), .I1(n3927), .S(n4897), .ZN(vectorData1[59])
         );
  MUX4ND0BWP U5856 ( .I0(\vrf/regTable[0][59] ), .I1(\vrf/regTable[1][59] ), 
        .I2(\vrf/regTable[2][59] ), .I3(\vrf/regTable[3][59] ), .S0(n4762), 
        .S1(n4832), .ZN(n3926) );
  MUX4ND0BWP U5857 ( .I0(\vrf/regTable[4][59] ), .I1(\vrf/regTable[5][59] ), 
        .I2(\vrf/regTable[6][59] ), .I3(\vrf/regTable[7][59] ), .S0(n4762), 
        .S1(n4832), .ZN(n3927) );
  MUX2ND0BWP U5858 ( .I0(n3928), .I1(n3929), .S(n4908), .ZN(vectorData1[187])
         );
  MUX4ND0BWP U5859 ( .I0(\vrf/regTable[0][187] ), .I1(\vrf/regTable[1][187] ), 
        .I2(\vrf/regTable[2][187] ), .I3(\vrf/regTable[3][187] ), .S0(n4784), 
        .S1(n4854), .ZN(n3928) );
  MUX4ND0BWP U5860 ( .I0(\vrf/regTable[4][187] ), .I1(\vrf/regTable[5][187] ), 
        .I2(\vrf/regTable[6][187] ), .I3(\vrf/regTable[7][187] ), .S0(n4784), 
        .S1(n4854), .ZN(n3929) );
  MUX2ND0BWP U5861 ( .I0(n3930), .I1(n3931), .S(n4903), .ZN(vectorData1[122])
         );
  MUX4ND0BWP U5862 ( .I0(\vrf/regTable[0][122] ), .I1(\vrf/regTable[1][122] ), 
        .I2(\vrf/regTable[2][122] ), .I3(\vrf/regTable[3][122] ), .S0(n4773), 
        .S1(n4843), .ZN(n3930) );
  MUX4ND0BWP U5863 ( .I0(\vrf/regTable[4][122] ), .I1(\vrf/regTable[5][122] ), 
        .I2(\vrf/regTable[6][122] ), .I3(\vrf/regTable[7][122] ), .S0(n4773), 
        .S1(n4843), .ZN(n3931) );
  MUX2ND0BWP U5864 ( .I0(n3932), .I1(n3933), .S(n4897), .ZN(vectorData1[58])
         );
  MUX4ND0BWP U5865 ( .I0(\vrf/regTable[0][58] ), .I1(\vrf/regTable[1][58] ), 
        .I2(\vrf/regTable[2][58] ), .I3(\vrf/regTable[3][58] ), .S0(n4762), 
        .S1(n4832), .ZN(n3932) );
  MUX4ND0BWP U5866 ( .I0(\vrf/regTable[4][58] ), .I1(\vrf/regTable[5][58] ), 
        .I2(\vrf/regTable[6][58] ), .I3(\vrf/regTable[7][58] ), .S0(n4762), 
        .S1(n4832), .ZN(n3933) );
  MUX2ND0BWP U5867 ( .I0(n3934), .I1(n3935), .S(n4908), .ZN(vectorData1[186])
         );
  MUX4ND0BWP U5868 ( .I0(\vrf/regTable[0][186] ), .I1(\vrf/regTable[1][186] ), 
        .I2(\vrf/regTable[2][186] ), .I3(\vrf/regTable[3][186] ), .S0(n4784), 
        .S1(n4854), .ZN(n3934) );
  MUX4ND0BWP U5869 ( .I0(\vrf/regTable[4][186] ), .I1(\vrf/regTable[5][186] ), 
        .I2(\vrf/regTable[6][186] ), .I3(\vrf/regTable[7][186] ), .S0(n4784), 
        .S1(n4854), .ZN(n3935) );
  MUX2ND0BWP U5870 ( .I0(n3936), .I1(n3937), .S(n4903), .ZN(vectorData1[121])
         );
  MUX4ND0BWP U5871 ( .I0(\vrf/regTable[0][121] ), .I1(\vrf/regTable[1][121] ), 
        .I2(\vrf/regTable[2][121] ), .I3(\vrf/regTable[3][121] ), .S0(n4773), 
        .S1(n4843), .ZN(n3936) );
  MUX4ND0BWP U5872 ( .I0(\vrf/regTable[4][121] ), .I1(\vrf/regTable[5][121] ), 
        .I2(\vrf/regTable[6][121] ), .I3(\vrf/regTable[7][121] ), .S0(n4773), 
        .S1(n4843), .ZN(n3937) );
  MUX2ND0BWP U5873 ( .I0(n3938), .I1(n3939), .S(n4897), .ZN(vectorData1[57])
         );
  MUX4ND0BWP U5874 ( .I0(\vrf/regTable[0][57] ), .I1(\vrf/regTable[1][57] ), 
        .I2(\vrf/regTable[2][57] ), .I3(\vrf/regTable[3][57] ), .S0(n4762), 
        .S1(n4832), .ZN(n3938) );
  MUX4ND0BWP U5875 ( .I0(\vrf/regTable[4][57] ), .I1(\vrf/regTable[5][57] ), 
        .I2(\vrf/regTable[6][57] ), .I3(\vrf/regTable[7][57] ), .S0(n4762), 
        .S1(n4832), .ZN(n3939) );
  MUX2ND0BWP U5876 ( .I0(n3940), .I1(n3941), .S(n4908), .ZN(vectorData1[185])
         );
  MUX4ND0BWP U5877 ( .I0(\vrf/regTable[0][185] ), .I1(\vrf/regTable[1][185] ), 
        .I2(\vrf/regTable[2][185] ), .I3(\vrf/regTable[3][185] ), .S0(n4783), 
        .S1(n4853), .ZN(n3940) );
  MUX4ND0BWP U5878 ( .I0(\vrf/regTable[4][185] ), .I1(\vrf/regTable[5][185] ), 
        .I2(\vrf/regTable[6][185] ), .I3(\vrf/regTable[7][185] ), .S0(n4783), 
        .S1(n4853), .ZN(n3941) );
  MUX2ND0BWP U5879 ( .I0(n3942), .I1(n3943), .S(n4903), .ZN(vectorData1[120])
         );
  MUX4ND0BWP U5880 ( .I0(\vrf/regTable[0][120] ), .I1(\vrf/regTable[1][120] ), 
        .I2(\vrf/regTable[2][120] ), .I3(\vrf/regTable[3][120] ), .S0(n4773), 
        .S1(n4843), .ZN(n3942) );
  MUX4ND0BWP U5881 ( .I0(\vrf/regTable[4][120] ), .I1(\vrf/regTable[5][120] ), 
        .I2(\vrf/regTable[6][120] ), .I3(\vrf/regTable[7][120] ), .S0(n4773), 
        .S1(n4843), .ZN(n3943) );
  MUX2ND0BWP U5882 ( .I0(n3944), .I1(n3945), .S(n4897), .ZN(vectorData1[56])
         );
  MUX4ND0BWP U5883 ( .I0(\vrf/regTable[0][56] ), .I1(\vrf/regTable[1][56] ), 
        .I2(\vrf/regTable[2][56] ), .I3(\vrf/regTable[3][56] ), .S0(n4762), 
        .S1(n4832), .ZN(n3944) );
  MUX4ND0BWP U5884 ( .I0(\vrf/regTable[4][56] ), .I1(\vrf/regTable[5][56] ), 
        .I2(\vrf/regTable[6][56] ), .I3(\vrf/regTable[7][56] ), .S0(n4762), 
        .S1(n4832), .ZN(n3945) );
  MUX2ND0BWP U5885 ( .I0(n3946), .I1(n3947), .S(n4908), .ZN(vectorData1[184])
         );
  MUX4ND0BWP U5886 ( .I0(\vrf/regTable[0][184] ), .I1(\vrf/regTable[1][184] ), 
        .I2(\vrf/regTable[2][184] ), .I3(\vrf/regTable[3][184] ), .S0(n4783), 
        .S1(n4853), .ZN(n3946) );
  MUX4ND0BWP U5887 ( .I0(\vrf/regTable[4][184] ), .I1(\vrf/regTable[5][184] ), 
        .I2(\vrf/regTable[6][184] ), .I3(\vrf/regTable[7][184] ), .S0(n4783), 
        .S1(n4853), .ZN(n3947) );
  MUX2ND0BWP U5888 ( .I0(n3948), .I1(n3949), .S(n4902), .ZN(vectorData1[113])
         );
  MUX4ND0BWP U5889 ( .I0(\vrf/regTable[0][113] ), .I1(\vrf/regTable[1][113] ), 
        .I2(\vrf/regTable[2][113] ), .I3(\vrf/regTable[3][113] ), .S0(n4771), 
        .S1(n4841), .ZN(n3948) );
  MUX4ND0BWP U5890 ( .I0(\vrf/regTable[4][113] ), .I1(\vrf/regTable[5][113] ), 
        .I2(\vrf/regTable[6][113] ), .I3(\vrf/regTable[7][113] ), .S0(n4771), 
        .S1(n4841), .ZN(n3949) );
  MUX2ND0BWP U5891 ( .I0(n3950), .I1(n3951), .S(n4897), .ZN(vectorData1[49])
         );
  MUX4ND0BWP U5892 ( .I0(\vrf/regTable[0][49] ), .I1(\vrf/regTable[1][49] ), 
        .I2(\vrf/regTable[2][49] ), .I3(\vrf/regTable[3][49] ), .S0(n4761), 
        .S1(n4831), .ZN(n3950) );
  MUX4ND0BWP U5893 ( .I0(\vrf/regTable[4][49] ), .I1(\vrf/regTable[5][49] ), 
        .I2(\vrf/regTable[6][49] ), .I3(\vrf/regTable[7][49] ), .S0(n4761), 
        .S1(n4831), .ZN(n3951) );
  MUX2ND0BWP U5894 ( .I0(n3952), .I1(n3953), .S(n4907), .ZN(vectorData1[177])
         );
  MUX4ND0BWP U5895 ( .I0(\vrf/regTable[0][177] ), .I1(\vrf/regTable[1][177] ), 
        .I2(\vrf/regTable[2][177] ), .I3(\vrf/regTable[3][177] ), .S0(n4782), 
        .S1(n4852), .ZN(n3952) );
  MUX4ND0BWP U5896 ( .I0(\vrf/regTable[4][177] ), .I1(\vrf/regTable[5][177] ), 
        .I2(\vrf/regTable[6][177] ), .I3(\vrf/regTable[7][177] ), .S0(n4782), 
        .S1(n4852), .ZN(n3953) );
  MUX2ND0BWP U5897 ( .I0(n3954), .I1(n3955), .S(n4902), .ZN(vectorData1[119])
         );
  MUX4ND0BWP U5898 ( .I0(\vrf/regTable[0][119] ), .I1(\vrf/regTable[1][119] ), 
        .I2(\vrf/regTable[2][119] ), .I3(\vrf/regTable[3][119] ), .S0(n4772), 
        .S1(n4842), .ZN(n3954) );
  MUX4ND0BWP U5899 ( .I0(\vrf/regTable[4][119] ), .I1(\vrf/regTable[5][119] ), 
        .I2(\vrf/regTable[6][119] ), .I3(\vrf/regTable[7][119] ), .S0(n4772), 
        .S1(n4842), .ZN(n3955) );
  MUX2ND0BWP U5900 ( .I0(n3956), .I1(n3957), .S(n4897), .ZN(vectorData1[55])
         );
  MUX4ND0BWP U5901 ( .I0(\vrf/regTable[0][55] ), .I1(\vrf/regTable[1][55] ), 
        .I2(\vrf/regTable[2][55] ), .I3(\vrf/regTable[3][55] ), .S0(n4762), 
        .S1(n4832), .ZN(n3956) );
  MUX4ND0BWP U5902 ( .I0(\vrf/regTable[4][55] ), .I1(\vrf/regTable[5][55] ), 
        .I2(\vrf/regTable[6][55] ), .I3(\vrf/regTable[7][55] ), .S0(n4762), 
        .S1(n4832), .ZN(n3957) );
  MUX2ND0BWP U5903 ( .I0(n3958), .I1(n3959), .S(n4908), .ZN(vectorData1[183])
         );
  MUX4ND0BWP U5904 ( .I0(\vrf/regTable[0][183] ), .I1(\vrf/regTable[1][183] ), 
        .I2(\vrf/regTable[2][183] ), .I3(\vrf/regTable[3][183] ), .S0(n4783), 
        .S1(n4853), .ZN(n3958) );
  MUX4ND0BWP U5905 ( .I0(\vrf/regTable[4][183] ), .I1(\vrf/regTable[5][183] ), 
        .I2(\vrf/regTable[6][183] ), .I3(\vrf/regTable[7][183] ), .S0(n4783), 
        .S1(n4853), .ZN(n3959) );
  MUX2ND0BWP U5906 ( .I0(n3960), .I1(n3961), .S(n4902), .ZN(vectorData1[118])
         );
  MUX4ND0BWP U5907 ( .I0(\vrf/regTable[0][118] ), .I1(\vrf/regTable[1][118] ), 
        .I2(\vrf/regTable[2][118] ), .I3(\vrf/regTable[3][118] ), .S0(n4772), 
        .S1(n4842), .ZN(n3960) );
  MUX4ND0BWP U5908 ( .I0(\vrf/regTable[4][118] ), .I1(\vrf/regTable[5][118] ), 
        .I2(\vrf/regTable[6][118] ), .I3(\vrf/regTable[7][118] ), .S0(n4772), 
        .S1(n4842), .ZN(n3961) );
  MUX2ND0BWP U5909 ( .I0(n3962), .I1(n3963), .S(n4897), .ZN(vectorData1[54])
         );
  MUX4ND0BWP U5910 ( .I0(\vrf/regTable[0][54] ), .I1(\vrf/regTable[1][54] ), 
        .I2(\vrf/regTable[2][54] ), .I3(\vrf/regTable[3][54] ), .S0(n4762), 
        .S1(n4832), .ZN(n3962) );
  MUX4ND0BWP U5911 ( .I0(\vrf/regTable[4][54] ), .I1(\vrf/regTable[5][54] ), 
        .I2(\vrf/regTable[6][54] ), .I3(\vrf/regTable[7][54] ), .S0(n4762), 
        .S1(n4832), .ZN(n3963) );
  MUX2ND0BWP U5912 ( .I0(n3964), .I1(n3965), .S(n4908), .ZN(vectorData1[182])
         );
  MUX4ND0BWP U5913 ( .I0(\vrf/regTable[0][182] ), .I1(\vrf/regTable[1][182] ), 
        .I2(\vrf/regTable[2][182] ), .I3(\vrf/regTable[3][182] ), .S0(n4783), 
        .S1(n4853), .ZN(n3964) );
  MUX4ND0BWP U5914 ( .I0(\vrf/regTable[4][182] ), .I1(\vrf/regTable[5][182] ), 
        .I2(\vrf/regTable[6][182] ), .I3(\vrf/regTable[7][182] ), .S0(n4783), 
        .S1(n4853), .ZN(n3965) );
  MUX2ND0BWP U5915 ( .I0(n3966), .I1(n3967), .S(n4902), .ZN(vectorData1[117])
         );
  MUX4ND0BWP U5916 ( .I0(\vrf/regTable[0][117] ), .I1(\vrf/regTable[1][117] ), 
        .I2(\vrf/regTable[2][117] ), .I3(\vrf/regTable[3][117] ), .S0(n4772), 
        .S1(n4842), .ZN(n3966) );
  MUX4ND0BWP U5917 ( .I0(\vrf/regTable[4][117] ), .I1(\vrf/regTable[5][117] ), 
        .I2(\vrf/regTable[6][117] ), .I3(\vrf/regTable[7][117] ), .S0(n4772), 
        .S1(n4842), .ZN(n3967) );
  MUX2ND0BWP U5918 ( .I0(n3968), .I1(n3969), .S(n4897), .ZN(vectorData1[53])
         );
  MUX4ND0BWP U5919 ( .I0(\vrf/regTable[0][53] ), .I1(\vrf/regTable[1][53] ), 
        .I2(\vrf/regTable[2][53] ), .I3(\vrf/regTable[3][53] ), .S0(n4761), 
        .S1(n4831), .ZN(n3968) );
  MUX4ND0BWP U5920 ( .I0(\vrf/regTable[4][53] ), .I1(\vrf/regTable[5][53] ), 
        .I2(\vrf/regTable[6][53] ), .I3(\vrf/regTable[7][53] ), .S0(n4761), 
        .S1(n4831), .ZN(n3969) );
  MUX2ND0BWP U5921 ( .I0(n3970), .I1(n3971), .S(n4908), .ZN(vectorData1[181])
         );
  MUX4ND0BWP U5922 ( .I0(\vrf/regTable[0][181] ), .I1(\vrf/regTable[1][181] ), 
        .I2(\vrf/regTable[2][181] ), .I3(\vrf/regTable[3][181] ), .S0(n4783), 
        .S1(n4853), .ZN(n3970) );
  MUX4ND0BWP U5923 ( .I0(\vrf/regTable[4][181] ), .I1(\vrf/regTable[5][181] ), 
        .I2(\vrf/regTable[6][181] ), .I3(\vrf/regTable[7][181] ), .S0(n4783), 
        .S1(n4853), .ZN(n3971) );
  MUX2ND0BWP U5924 ( .I0(n3972), .I1(n3973), .S(n4902), .ZN(vectorData1[114])
         );
  MUX4ND0BWP U5925 ( .I0(\vrf/regTable[0][114] ), .I1(\vrf/regTable[1][114] ), 
        .I2(\vrf/regTable[2][114] ), .I3(\vrf/regTable[3][114] ), .S0(n4772), 
        .S1(n4842), .ZN(n3972) );
  MUX4ND0BWP U5926 ( .I0(\vrf/regTable[4][114] ), .I1(\vrf/regTable[5][114] ), 
        .I2(\vrf/regTable[6][114] ), .I3(\vrf/regTable[7][114] ), .S0(n4772), 
        .S1(n4842), .ZN(n3973) );
  MUX2ND0BWP U5927 ( .I0(n3974), .I1(n3975), .S(n4897), .ZN(vectorData1[50])
         );
  MUX4ND0BWP U5928 ( .I0(\vrf/regTable[0][50] ), .I1(\vrf/regTable[1][50] ), 
        .I2(\vrf/regTable[2][50] ), .I3(\vrf/regTable[3][50] ), .S0(n4761), 
        .S1(n4831), .ZN(n3974) );
  MUX4ND0BWP U5929 ( .I0(\vrf/regTable[4][50] ), .I1(\vrf/regTable[5][50] ), 
        .I2(\vrf/regTable[6][50] ), .I3(\vrf/regTable[7][50] ), .S0(n4761), 
        .S1(n4831), .ZN(n3975) );
  MUX2ND0BWP U5930 ( .I0(n3976), .I1(n3977), .S(n4907), .ZN(vectorData1[178])
         );
  MUX4ND0BWP U5931 ( .I0(\vrf/regTable[0][178] ), .I1(\vrf/regTable[1][178] ), 
        .I2(\vrf/regTable[2][178] ), .I3(\vrf/regTable[3][178] ), .S0(n4782), 
        .S1(n4852), .ZN(n3976) );
  MUX4ND0BWP U5932 ( .I0(\vrf/regTable[4][178] ), .I1(\vrf/regTable[5][178] ), 
        .I2(\vrf/regTable[6][178] ), .I3(\vrf/regTable[7][178] ), .S0(n4782), 
        .S1(n4852), .ZN(n3977) );
  MUX2ND0BWP U5933 ( .I0(n3978), .I1(n3979), .S(n4902), .ZN(vectorData1[115])
         );
  MUX4ND0BWP U5934 ( .I0(\vrf/regTable[0][115] ), .I1(\vrf/regTable[1][115] ), 
        .I2(\vrf/regTable[2][115] ), .I3(\vrf/regTable[3][115] ), .S0(n4772), 
        .S1(n4842), .ZN(n3978) );
  MUX4ND0BWP U5935 ( .I0(\vrf/regTable[4][115] ), .I1(\vrf/regTable[5][115] ), 
        .I2(\vrf/regTable[6][115] ), .I3(\vrf/regTable[7][115] ), .S0(n4772), 
        .S1(n4842), .ZN(n3979) );
  MUX2ND0BWP U5936 ( .I0(n3980), .I1(n3981), .S(n4897), .ZN(vectorData1[51])
         );
  MUX4ND0BWP U5937 ( .I0(\vrf/regTable[0][51] ), .I1(\vrf/regTable[1][51] ), 
        .I2(\vrf/regTable[2][51] ), .I3(\vrf/regTable[3][51] ), .S0(n4761), 
        .S1(n4831), .ZN(n3980) );
  MUX4ND0BWP U5938 ( .I0(\vrf/regTable[4][51] ), .I1(\vrf/regTable[5][51] ), 
        .I2(\vrf/regTable[6][51] ), .I3(\vrf/regTable[7][51] ), .S0(n4761), 
        .S1(n4831), .ZN(n3981) );
  MUX2ND0BWP U5939 ( .I0(n3982), .I1(n3983), .S(n4907), .ZN(vectorData1[179])
         );
  MUX4ND0BWP U5940 ( .I0(\vrf/regTable[0][179] ), .I1(\vrf/regTable[1][179] ), 
        .I2(\vrf/regTable[2][179] ), .I3(\vrf/regTable[3][179] ), .S0(n4782), 
        .S1(n4852), .ZN(n3982) );
  MUX4ND0BWP U5941 ( .I0(\vrf/regTable[4][179] ), .I1(\vrf/regTable[5][179] ), 
        .I2(\vrf/regTable[6][179] ), .I3(\vrf/regTable[7][179] ), .S0(n4782), 
        .S1(n4852), .ZN(n3983) );
  MUX2ND0BWP U5942 ( .I0(n3984), .I1(n3985), .S(n4902), .ZN(vectorData1[116])
         );
  MUX4ND0BWP U5943 ( .I0(\vrf/regTable[0][116] ), .I1(\vrf/regTable[1][116] ), 
        .I2(\vrf/regTable[2][116] ), .I3(\vrf/regTable[3][116] ), .S0(n4772), 
        .S1(n4842), .ZN(n3984) );
  MUX4ND0BWP U5944 ( .I0(\vrf/regTable[4][116] ), .I1(\vrf/regTable[5][116] ), 
        .I2(\vrf/regTable[6][116] ), .I3(\vrf/regTable[7][116] ), .S0(n4772), 
        .S1(n4842), .ZN(n3985) );
  MUX2ND0BWP U5945 ( .I0(n3986), .I1(n3987), .S(n4897), .ZN(vectorData1[52])
         );
  MUX4ND0BWP U5946 ( .I0(\vrf/regTable[0][52] ), .I1(\vrf/regTable[1][52] ), 
        .I2(\vrf/regTable[2][52] ), .I3(\vrf/regTable[3][52] ), .S0(n4761), 
        .S1(n4831), .ZN(n3986) );
  MUX4ND0BWP U5947 ( .I0(\vrf/regTable[4][52] ), .I1(\vrf/regTable[5][52] ), 
        .I2(\vrf/regTable[6][52] ), .I3(\vrf/regTable[7][52] ), .S0(n4761), 
        .S1(n4831), .ZN(n3987) );
  MUX2ND0BWP U5948 ( .I0(n3988), .I1(n3989), .S(n4908), .ZN(vectorData1[180])
         );
  MUX4ND0BWP U5949 ( .I0(\vrf/regTable[0][180] ), .I1(\vrf/regTable[1][180] ), 
        .I2(\vrf/regTable[2][180] ), .I3(\vrf/regTable[3][180] ), .S0(n4783), 
        .S1(n4853), .ZN(n3988) );
  MUX4ND0BWP U5950 ( .I0(\vrf/regTable[4][180] ), .I1(\vrf/regTable[5][180] ), 
        .I2(\vrf/regTable[6][180] ), .I3(\vrf/regTable[7][180] ), .S0(n4783), 
        .S1(n4853), .ZN(n3989) );
  MUX2ND0BWP U5951 ( .I0(n3990), .I1(n3991), .S(n4901), .ZN(vectorData1[96])
         );
  MUX4ND0BWP U5952 ( .I0(\vrf/regTable[0][96] ), .I1(\vrf/regTable[1][96] ), 
        .I2(\vrf/regTable[2][96] ), .I3(\vrf/regTable[3][96] ), .S0(n4769), 
        .S1(n4839), .ZN(n3990) );
  MUX4ND0BWP U5953 ( .I0(\vrf/regTable[4][96] ), .I1(\vrf/regTable[5][96] ), 
        .I2(\vrf/regTable[6][96] ), .I3(\vrf/regTable[7][96] ), .S0(n4769), 
        .S1(n4839), .ZN(n3991) );
  MUX2ND0BWP U5954 ( .I0(n3992), .I1(n3993), .S(n4895), .ZN(vectorData1[32])
         );
  MUX4ND0BWP U5955 ( .I0(\vrf/regTable[0][32] ), .I1(\vrf/regTable[1][32] ), 
        .I2(\vrf/regTable[2][32] ), .I3(\vrf/regTable[3][32] ), .S0(n4758), 
        .S1(n4828), .ZN(n3992) );
  MUX4ND0BWP U5956 ( .I0(\vrf/regTable[4][32] ), .I1(\vrf/regTable[5][32] ), 
        .I2(\vrf/regTable[6][32] ), .I3(\vrf/regTable[7][32] ), .S0(n4758), 
        .S1(n4828), .ZN(n3993) );
  MUX2ND0BWP U5957 ( .I0(n3994), .I1(n3995), .S(n4906), .ZN(vectorData1[160])
         );
  MUX4ND0BWP U5958 ( .I0(\vrf/regTable[0][160] ), .I1(\vrf/regTable[1][160] ), 
        .I2(\vrf/regTable[2][160] ), .I3(\vrf/regTable[3][160] ), .S0(n4779), 
        .S1(n4849), .ZN(n3994) );
  MUX4ND0BWP U5959 ( .I0(\vrf/regTable[4][160] ), .I1(\vrf/regTable[5][160] ), 
        .I2(\vrf/regTable[6][160] ), .I3(\vrf/regTable[7][160] ), .S0(n4779), 
        .S1(n4849), .ZN(n3995) );
  MUX2ND0BWP U5960 ( .I0(n3996), .I1(n3997), .S(n4902), .ZN(vectorData1[111])
         );
  MUX4ND0BWP U5961 ( .I0(\vrf/regTable[0][111] ), .I1(\vrf/regTable[1][111] ), 
        .I2(\vrf/regTable[2][111] ), .I3(\vrf/regTable[3][111] ), .S0(n4771), 
        .S1(n4841), .ZN(n3996) );
  MUX4ND0BWP U5962 ( .I0(\vrf/regTable[4][111] ), .I1(\vrf/regTable[5][111] ), 
        .I2(\vrf/regTable[6][111] ), .I3(\vrf/regTable[7][111] ), .S0(n4771), 
        .S1(n4841), .ZN(n3997) );
  MUX2ND0BWP U5963 ( .I0(n3998), .I1(n3999), .S(n4896), .ZN(vectorData1[47])
         );
  MUX4ND0BWP U5964 ( .I0(\vrf/regTable[0][47] ), .I1(\vrf/regTable[1][47] ), 
        .I2(\vrf/regTable[2][47] ), .I3(\vrf/regTable[3][47] ), .S0(n4760), 
        .S1(n4830), .ZN(n3998) );
  MUX4ND0BWP U5965 ( .I0(\vrf/regTable[4][47] ), .I1(\vrf/regTable[5][47] ), 
        .I2(\vrf/regTable[6][47] ), .I3(\vrf/regTable[7][47] ), .S0(n4760), 
        .S1(n4830), .ZN(n3999) );
  MUX2ND0BWP U5966 ( .I0(n4000), .I1(n4001), .S(n4907), .ZN(vectorData1[175])
         );
  MUX4ND0BWP U5967 ( .I0(\vrf/regTable[0][175] ), .I1(\vrf/regTable[1][175] ), 
        .I2(\vrf/regTable[2][175] ), .I3(\vrf/regTable[3][175] ), .S0(n4782), 
        .S1(n4852), .ZN(n4000) );
  MUX4ND0BWP U5968 ( .I0(\vrf/regTable[4][175] ), .I1(\vrf/regTable[5][175] ), 
        .I2(\vrf/regTable[6][175] ), .I3(\vrf/regTable[7][175] ), .S0(n4782), 
        .S1(n4852), .ZN(n4001) );
  MUX2ND0BWP U5969 ( .I0(n4002), .I1(n4003), .S(n4902), .ZN(vectorData1[110])
         );
  MUX4ND0BWP U5970 ( .I0(\vrf/regTable[0][110] ), .I1(\vrf/regTable[1][110] ), 
        .I2(\vrf/regTable[2][110] ), .I3(\vrf/regTable[3][110] ), .S0(n4771), 
        .S1(n4841), .ZN(n4002) );
  MUX4ND0BWP U5971 ( .I0(\vrf/regTable[4][110] ), .I1(\vrf/regTable[5][110] ), 
        .I2(\vrf/regTable[6][110] ), .I3(\vrf/regTable[7][110] ), .S0(n4771), 
        .S1(n4841), .ZN(n4003) );
  MUX2ND0BWP U5972 ( .I0(n4004), .I1(n4005), .S(n4896), .ZN(vectorData1[46])
         );
  MUX4ND0BWP U5973 ( .I0(\vrf/regTable[0][46] ), .I1(\vrf/regTable[1][46] ), 
        .I2(\vrf/regTable[2][46] ), .I3(\vrf/regTable[3][46] ), .S0(n4760), 
        .S1(n4830), .ZN(n4004) );
  MUX4ND0BWP U5974 ( .I0(\vrf/regTable[4][46] ), .I1(\vrf/regTable[5][46] ), 
        .I2(\vrf/regTable[6][46] ), .I3(\vrf/regTable[7][46] ), .S0(n4760), 
        .S1(n4830), .ZN(n4005) );
  MUX2ND0BWP U5975 ( .I0(n4006), .I1(n4007), .S(n4907), .ZN(vectorData1[174])
         );
  MUX4ND0BWP U5976 ( .I0(\vrf/regTable[0][174] ), .I1(\vrf/regTable[1][174] ), 
        .I2(\vrf/regTable[2][174] ), .I3(\vrf/regTable[3][174] ), .S0(n4782), 
        .S1(n4852), .ZN(n4006) );
  MUX4ND0BWP U5977 ( .I0(\vrf/regTable[4][174] ), .I1(\vrf/regTable[5][174] ), 
        .I2(\vrf/regTable[6][174] ), .I3(\vrf/regTable[7][174] ), .S0(n4782), 
        .S1(n4852), .ZN(n4007) );
  MUX2ND0BWP U5978 ( .I0(n4008), .I1(n4009), .S(n4902), .ZN(vectorData1[109])
         );
  MUX4ND0BWP U5979 ( .I0(\vrf/regTable[0][109] ), .I1(\vrf/regTable[1][109] ), 
        .I2(\vrf/regTable[2][109] ), .I3(\vrf/regTable[3][109] ), .S0(n4771), 
        .S1(n4841), .ZN(n4008) );
  MUX4ND0BWP U5980 ( .I0(\vrf/regTable[4][109] ), .I1(\vrf/regTable[5][109] ), 
        .I2(\vrf/regTable[6][109] ), .I3(\vrf/regTable[7][109] ), .S0(n4771), 
        .S1(n4841), .ZN(n4009) );
  MUX2ND0BWP U5981 ( .I0(n4010), .I1(n4011), .S(n4896), .ZN(vectorData1[45])
         );
  MUX4ND0BWP U5982 ( .I0(\vrf/regTable[0][45] ), .I1(\vrf/regTable[1][45] ), 
        .I2(\vrf/regTable[2][45] ), .I3(\vrf/regTable[3][45] ), .S0(n4760), 
        .S1(n4830), .ZN(n4010) );
  MUX4ND0BWP U5983 ( .I0(\vrf/regTable[4][45] ), .I1(\vrf/regTable[5][45] ), 
        .I2(\vrf/regTable[6][45] ), .I3(\vrf/regTable[7][45] ), .S0(n4760), 
        .S1(n4830), .ZN(n4011) );
  MUX2ND0BWP U5984 ( .I0(n4012), .I1(n4013), .S(n4907), .ZN(vectorData1[173])
         );
  MUX4ND0BWP U5985 ( .I0(\vrf/regTable[0][173] ), .I1(\vrf/regTable[1][173] ), 
        .I2(\vrf/regTable[2][173] ), .I3(\vrf/regTable[3][173] ), .S0(n4781), 
        .S1(n4851), .ZN(n4012) );
  MUX4ND0BWP U5986 ( .I0(\vrf/regTable[4][173] ), .I1(\vrf/regTable[5][173] ), 
        .I2(\vrf/regTable[6][173] ), .I3(\vrf/regTable[7][173] ), .S0(n4781), 
        .S1(n4851), .ZN(n4013) );
  MUX2ND0BWP U5987 ( .I0(n4014), .I1(n4015), .S(n4902), .ZN(vectorData1[108])
         );
  MUX4ND0BWP U5988 ( .I0(\vrf/regTable[0][108] ), .I1(\vrf/regTable[1][108] ), 
        .I2(\vrf/regTable[2][108] ), .I3(\vrf/regTable[3][108] ), .S0(n4771), 
        .S1(n4841), .ZN(n4014) );
  MUX4ND0BWP U5989 ( .I0(\vrf/regTable[4][108] ), .I1(\vrf/regTable[5][108] ), 
        .I2(\vrf/regTable[6][108] ), .I3(\vrf/regTable[7][108] ), .S0(n4771), 
        .S1(n4841), .ZN(n4015) );
  MUX2ND0BWP U5990 ( .I0(n4016), .I1(n4017), .S(n4896), .ZN(vectorData1[44])
         );
  MUX4ND0BWP U5991 ( .I0(\vrf/regTable[0][44] ), .I1(\vrf/regTable[1][44] ), 
        .I2(\vrf/regTable[2][44] ), .I3(\vrf/regTable[3][44] ), .S0(n4760), 
        .S1(n4830), .ZN(n4016) );
  MUX4ND0BWP U5992 ( .I0(\vrf/regTable[4][44] ), .I1(\vrf/regTable[5][44] ), 
        .I2(\vrf/regTable[6][44] ), .I3(\vrf/regTable[7][44] ), .S0(n4760), 
        .S1(n4830), .ZN(n4017) );
  MUX2ND0BWP U5993 ( .I0(n4018), .I1(n4019), .S(n4907), .ZN(vectorData1[172])
         );
  MUX4ND0BWP U5994 ( .I0(\vrf/regTable[0][172] ), .I1(\vrf/regTable[1][172] ), 
        .I2(\vrf/regTable[2][172] ), .I3(\vrf/regTable[3][172] ), .S0(n4781), 
        .S1(n4851), .ZN(n4018) );
  MUX4ND0BWP U5995 ( .I0(\vrf/regTable[4][172] ), .I1(\vrf/regTable[5][172] ), 
        .I2(\vrf/regTable[6][172] ), .I3(\vrf/regTable[7][172] ), .S0(n4781), 
        .S1(n4851), .ZN(n4019) );
  MUX2ND0BWP U5996 ( .I0(n4020), .I1(n4021), .S(n4901), .ZN(vectorData1[107])
         );
  MUX4ND0BWP U5997 ( .I0(\vrf/regTable[0][107] ), .I1(\vrf/regTable[1][107] ), 
        .I2(\vrf/regTable[2][107] ), .I3(\vrf/regTable[3][107] ), .S0(n4770), 
        .S1(n4840), .ZN(n4020) );
  MUX4ND0BWP U5998 ( .I0(\vrf/regTable[4][107] ), .I1(\vrf/regTable[5][107] ), 
        .I2(\vrf/regTable[6][107] ), .I3(\vrf/regTable[7][107] ), .S0(n4770), 
        .S1(n4840), .ZN(n4021) );
  MUX2ND0BWP U5999 ( .I0(n4022), .I1(n4023), .S(n4896), .ZN(vectorData1[43])
         );
  MUX4ND0BWP U6000 ( .I0(\vrf/regTable[0][43] ), .I1(\vrf/regTable[1][43] ), 
        .I2(\vrf/regTable[2][43] ), .I3(\vrf/regTable[3][43] ), .S0(n4760), 
        .S1(n4830), .ZN(n4022) );
  MUX4ND0BWP U6001 ( .I0(\vrf/regTable[4][43] ), .I1(\vrf/regTable[5][43] ), 
        .I2(\vrf/regTable[6][43] ), .I3(\vrf/regTable[7][43] ), .S0(n4760), 
        .S1(n4830), .ZN(n4023) );
  MUX2ND0BWP U6002 ( .I0(n4024), .I1(n4025), .S(n4907), .ZN(vectorData1[171])
         );
  MUX4ND0BWP U6003 ( .I0(\vrf/regTable[0][171] ), .I1(\vrf/regTable[1][171] ), 
        .I2(\vrf/regTable[2][171] ), .I3(\vrf/regTable[3][171] ), .S0(n4781), 
        .S1(n4851), .ZN(n4024) );
  MUX4ND0BWP U6004 ( .I0(\vrf/regTable[4][171] ), .I1(\vrf/regTable[5][171] ), 
        .I2(\vrf/regTable[6][171] ), .I3(\vrf/regTable[7][171] ), .S0(n4781), 
        .S1(n4851), .ZN(n4025) );
  MUX2ND0BWP U6005 ( .I0(n4026), .I1(n4027), .S(n4901), .ZN(vectorData1[106])
         );
  MUX4ND0BWP U6006 ( .I0(\vrf/regTable[0][106] ), .I1(\vrf/regTable[1][106] ), 
        .I2(\vrf/regTable[2][106] ), .I3(\vrf/regTable[3][106] ), .S0(n4770), 
        .S1(n4840), .ZN(n4026) );
  MUX4ND0BWP U6007 ( .I0(\vrf/regTable[4][106] ), .I1(\vrf/regTable[5][106] ), 
        .I2(\vrf/regTable[6][106] ), .I3(\vrf/regTable[7][106] ), .S0(n4770), 
        .S1(n4840), .ZN(n4027) );
  MUX2ND0BWP U6008 ( .I0(n4028), .I1(n4029), .S(n4896), .ZN(vectorData1[42])
         );
  MUX4ND0BWP U6009 ( .I0(\vrf/regTable[0][42] ), .I1(\vrf/regTable[1][42] ), 
        .I2(\vrf/regTable[2][42] ), .I3(\vrf/regTable[3][42] ), .S0(n4760), 
        .S1(n4830), .ZN(n4028) );
  MUX4ND0BWP U6010 ( .I0(\vrf/regTable[4][42] ), .I1(\vrf/regTable[5][42] ), 
        .I2(\vrf/regTable[6][42] ), .I3(\vrf/regTable[7][42] ), .S0(n4760), 
        .S1(n4830), .ZN(n4029) );
  MUX2ND0BWP U6011 ( .I0(n4030), .I1(n4031), .S(n4907), .ZN(vectorData1[170])
         );
  MUX4ND0BWP U6012 ( .I0(\vrf/regTable[0][170] ), .I1(\vrf/regTable[1][170] ), 
        .I2(\vrf/regTable[2][170] ), .I3(\vrf/regTable[3][170] ), .S0(n4781), 
        .S1(n4851), .ZN(n4030) );
  MUX4ND0BWP U6013 ( .I0(\vrf/regTable[4][170] ), .I1(\vrf/regTable[5][170] ), 
        .I2(\vrf/regTable[6][170] ), .I3(\vrf/regTable[7][170] ), .S0(n4781), 
        .S1(n4851), .ZN(n4031) );
  MUX2ND0BWP U6014 ( .I0(n4032), .I1(n4033), .S(n4901), .ZN(vectorData1[105])
         );
  MUX4ND0BWP U6015 ( .I0(\vrf/regTable[0][105] ), .I1(\vrf/regTable[1][105] ), 
        .I2(\vrf/regTable[2][105] ), .I3(\vrf/regTable[3][105] ), .S0(n4770), 
        .S1(n4840), .ZN(n4032) );
  MUX4ND0BWP U6016 ( .I0(\vrf/regTable[4][105] ), .I1(\vrf/regTable[5][105] ), 
        .I2(\vrf/regTable[6][105] ), .I3(\vrf/regTable[7][105] ), .S0(n4770), 
        .S1(n4840), .ZN(n4033) );
  MUX2ND0BWP U6017 ( .I0(n4034), .I1(n4035), .S(n4896), .ZN(vectorData1[41])
         );
  MUX4ND0BWP U6018 ( .I0(\vrf/regTable[0][41] ), .I1(\vrf/regTable[1][41] ), 
        .I2(\vrf/regTable[2][41] ), .I3(\vrf/regTable[3][41] ), .S0(n4759), 
        .S1(n4829), .ZN(n4034) );
  MUX4ND0BWP U6019 ( .I0(\vrf/regTable[4][41] ), .I1(\vrf/regTable[5][41] ), 
        .I2(\vrf/regTable[6][41] ), .I3(\vrf/regTable[7][41] ), .S0(n4759), 
        .S1(n4829), .ZN(n4035) );
  MUX2ND0BWP U6020 ( .I0(n4036), .I1(n4037), .S(n4907), .ZN(vectorData1[169])
         );
  MUX4ND0BWP U6021 ( .I0(\vrf/regTable[0][169] ), .I1(\vrf/regTable[1][169] ), 
        .I2(\vrf/regTable[2][169] ), .I3(\vrf/regTable[3][169] ), .S0(n4781), 
        .S1(n4851), .ZN(n4036) );
  MUX4ND0BWP U6022 ( .I0(\vrf/regTable[4][169] ), .I1(\vrf/regTable[5][169] ), 
        .I2(\vrf/regTable[6][169] ), .I3(\vrf/regTable[7][169] ), .S0(n4781), 
        .S1(n4851), .ZN(n4037) );
  MUX2ND0BWP U6023 ( .I0(n4038), .I1(n4039), .S(n4901), .ZN(vectorData1[104])
         );
  MUX4ND0BWP U6024 ( .I0(\vrf/regTable[0][104] ), .I1(\vrf/regTable[1][104] ), 
        .I2(\vrf/regTable[2][104] ), .I3(\vrf/regTable[3][104] ), .S0(n4770), 
        .S1(n4840), .ZN(n4038) );
  MUX4ND0BWP U6025 ( .I0(\vrf/regTable[4][104] ), .I1(\vrf/regTable[5][104] ), 
        .I2(\vrf/regTable[6][104] ), .I3(\vrf/regTable[7][104] ), .S0(n4770), 
        .S1(n4840), .ZN(n4039) );
  MUX2ND0BWP U6026 ( .I0(n4040), .I1(n4041), .S(n4896), .ZN(vectorData1[40])
         );
  MUX4ND0BWP U6027 ( .I0(\vrf/regTable[0][40] ), .I1(\vrf/regTable[1][40] ), 
        .I2(\vrf/regTable[2][40] ), .I3(\vrf/regTable[3][40] ), .S0(n4759), 
        .S1(n4829), .ZN(n4040) );
  MUX4ND0BWP U6028 ( .I0(\vrf/regTable[4][40] ), .I1(\vrf/regTable[5][40] ), 
        .I2(\vrf/regTable[6][40] ), .I3(\vrf/regTable[7][40] ), .S0(n4759), 
        .S1(n4829), .ZN(n4041) );
  MUX2ND0BWP U6029 ( .I0(n4042), .I1(n4043), .S(n4907), .ZN(vectorData1[168])
         );
  MUX4ND0BWP U6030 ( .I0(\vrf/regTable[0][168] ), .I1(\vrf/regTable[1][168] ), 
        .I2(\vrf/regTable[2][168] ), .I3(\vrf/regTable[3][168] ), .S0(n4781), 
        .S1(n4851), .ZN(n4042) );
  MUX4ND0BWP U6031 ( .I0(\vrf/regTable[4][168] ), .I1(\vrf/regTable[5][168] ), 
        .I2(\vrf/regTable[6][168] ), .I3(\vrf/regTable[7][168] ), .S0(n4781), 
        .S1(n4851), .ZN(n4043) );
  MUX2ND0BWP U6032 ( .I0(n4044), .I1(n4045), .S(n4901), .ZN(vectorData1[97])
         );
  MUX4ND0BWP U6033 ( .I0(\vrf/regTable[0][97] ), .I1(\vrf/regTable[1][97] ), 
        .I2(\vrf/regTable[2][97] ), .I3(\vrf/regTable[3][97] ), .S0(n4769), 
        .S1(n4839), .ZN(n4044) );
  MUX4ND0BWP U6034 ( .I0(\vrf/regTable[4][97] ), .I1(\vrf/regTable[5][97] ), 
        .I2(\vrf/regTable[6][97] ), .I3(\vrf/regTable[7][97] ), .S0(n4769), 
        .S1(n4839), .ZN(n4045) );
  MUX2ND0BWP U6035 ( .I0(n4046), .I1(n4047), .S(n4895), .ZN(vectorData1[33])
         );
  MUX4ND0BWP U6036 ( .I0(\vrf/regTable[0][33] ), .I1(\vrf/regTable[1][33] ), 
        .I2(\vrf/regTable[2][33] ), .I3(\vrf/regTable[3][33] ), .S0(n4758), 
        .S1(n4828), .ZN(n4046) );
  MUX4ND0BWP U6037 ( .I0(\vrf/regTable[4][33] ), .I1(\vrf/regTable[5][33] ), 
        .I2(\vrf/regTable[6][33] ), .I3(\vrf/regTable[7][33] ), .S0(n4758), 
        .S1(n4828), .ZN(n4047) );
  MUX2ND0BWP U6038 ( .I0(n4048), .I1(n4049), .S(n4906), .ZN(vectorData1[161])
         );
  MUX4ND0BWP U6039 ( .I0(\vrf/regTable[0][161] ), .I1(\vrf/regTable[1][161] ), 
        .I2(\vrf/regTable[2][161] ), .I3(\vrf/regTable[3][161] ), .S0(n4779), 
        .S1(n4849), .ZN(n4048) );
  MUX4ND0BWP U6040 ( .I0(\vrf/regTable[4][161] ), .I1(\vrf/regTable[5][161] ), 
        .I2(\vrf/regTable[6][161] ), .I3(\vrf/regTable[7][161] ), .S0(n4779), 
        .S1(n4849), .ZN(n4049) );
  MUX2ND0BWP U6041 ( .I0(n4050), .I1(n4051), .S(n4901), .ZN(vectorData1[103])
         );
  MUX4ND0BWP U6042 ( .I0(\vrf/regTable[0][103] ), .I1(\vrf/regTable[1][103] ), 
        .I2(\vrf/regTable[2][103] ), .I3(\vrf/regTable[3][103] ), .S0(n4770), 
        .S1(n4840), .ZN(n4050) );
  MUX4ND0BWP U6043 ( .I0(\vrf/regTable[4][103] ), .I1(\vrf/regTable[5][103] ), 
        .I2(\vrf/regTable[6][103] ), .I3(\vrf/regTable[7][103] ), .S0(n4770), 
        .S1(n4840), .ZN(n4051) );
  MUX2ND0BWP U6044 ( .I0(n4052), .I1(n4053), .S(n4896), .ZN(vectorData1[39])
         );
  MUX4ND0BWP U6045 ( .I0(\vrf/regTable[0][39] ), .I1(\vrf/regTable[1][39] ), 
        .I2(\vrf/regTable[2][39] ), .I3(\vrf/regTable[3][39] ), .S0(n4759), 
        .S1(n4829), .ZN(n4052) );
  MUX4ND0BWP U6046 ( .I0(\vrf/regTable[4][39] ), .I1(\vrf/regTable[5][39] ), 
        .I2(\vrf/regTable[6][39] ), .I3(\vrf/regTable[7][39] ), .S0(n4759), 
        .S1(n4829), .ZN(n4053) );
  MUX2ND0BWP U6047 ( .I0(n4054), .I1(n4055), .S(n4906), .ZN(vectorData1[167])
         );
  MUX4ND0BWP U6048 ( .I0(\vrf/regTable[0][167] ), .I1(\vrf/regTable[1][167] ), 
        .I2(\vrf/regTable[2][167] ), .I3(\vrf/regTable[3][167] ), .S0(n4780), 
        .S1(n4850), .ZN(n4054) );
  MUX4ND0BWP U6049 ( .I0(\vrf/regTable[4][167] ), .I1(\vrf/regTable[5][167] ), 
        .I2(\vrf/regTable[6][167] ), .I3(\vrf/regTable[7][167] ), .S0(n4780), 
        .S1(n4850), .ZN(n4055) );
  MUX2ND0BWP U6050 ( .I0(n4056), .I1(n4057), .S(n4901), .ZN(vectorData1[102])
         );
  MUX4ND0BWP U6051 ( .I0(\vrf/regTable[0][102] ), .I1(\vrf/regTable[1][102] ), 
        .I2(\vrf/regTable[2][102] ), .I3(\vrf/regTable[3][102] ), .S0(n4770), 
        .S1(n4840), .ZN(n4056) );
  MUX4ND0BWP U6052 ( .I0(\vrf/regTable[4][102] ), .I1(\vrf/regTable[5][102] ), 
        .I2(\vrf/regTable[6][102] ), .I3(\vrf/regTable[7][102] ), .S0(n4770), 
        .S1(n4840), .ZN(n4057) );
  MUX2ND0BWP U6053 ( .I0(n4058), .I1(n4059), .S(n4896), .ZN(vectorData1[38])
         );
  MUX4ND0BWP U6054 ( .I0(\vrf/regTable[0][38] ), .I1(\vrf/regTable[1][38] ), 
        .I2(\vrf/regTable[2][38] ), .I3(\vrf/regTable[3][38] ), .S0(n4759), 
        .S1(n4829), .ZN(n4058) );
  MUX4ND0BWP U6055 ( .I0(\vrf/regTable[4][38] ), .I1(\vrf/regTable[5][38] ), 
        .I2(\vrf/regTable[6][38] ), .I3(\vrf/regTable[7][38] ), .S0(n4759), 
        .S1(n4829), .ZN(n4059) );
  MUX2ND0BWP U6056 ( .I0(n4060), .I1(n4061), .S(n4906), .ZN(vectorData1[166])
         );
  MUX4ND0BWP U6057 ( .I0(\vrf/regTable[0][166] ), .I1(\vrf/regTable[1][166] ), 
        .I2(\vrf/regTable[2][166] ), .I3(\vrf/regTable[3][166] ), .S0(n4780), 
        .S1(n4850), .ZN(n4060) );
  MUX4ND0BWP U6058 ( .I0(\vrf/regTable[4][166] ), .I1(\vrf/regTable[5][166] ), 
        .I2(\vrf/regTable[6][166] ), .I3(\vrf/regTable[7][166] ), .S0(n4780), 
        .S1(n4850), .ZN(n4061) );
  MUX2ND0BWP U6059 ( .I0(n4062), .I1(n4063), .S(n4901), .ZN(vectorData1[101])
         );
  MUX4ND0BWP U6060 ( .I0(\vrf/regTable[0][101] ), .I1(\vrf/regTable[1][101] ), 
        .I2(\vrf/regTable[2][101] ), .I3(\vrf/regTable[3][101] ), .S0(n4769), 
        .S1(n4839), .ZN(n4062) );
  MUX4ND0BWP U6061 ( .I0(\vrf/regTable[4][101] ), .I1(\vrf/regTable[5][101] ), 
        .I2(\vrf/regTable[6][101] ), .I3(\vrf/regTable[7][101] ), .S0(n4769), 
        .S1(n4839), .ZN(n4063) );
  MUX2ND0BWP U6062 ( .I0(n4064), .I1(n4065), .S(n4896), .ZN(vectorData1[37])
         );
  MUX4ND0BWP U6063 ( .I0(\vrf/regTable[0][37] ), .I1(\vrf/regTable[1][37] ), 
        .I2(\vrf/regTable[2][37] ), .I3(\vrf/regTable[3][37] ), .S0(n4759), 
        .S1(n4829), .ZN(n4064) );
  MUX4ND0BWP U6064 ( .I0(\vrf/regTable[4][37] ), .I1(\vrf/regTable[5][37] ), 
        .I2(\vrf/regTable[6][37] ), .I3(\vrf/regTable[7][37] ), .S0(n4759), 
        .S1(n4829), .ZN(n4065) );
  MUX2ND0BWP U6065 ( .I0(n4066), .I1(n4067), .S(n4906), .ZN(vectorData1[165])
         );
  MUX4ND0BWP U6066 ( .I0(\vrf/regTable[0][165] ), .I1(\vrf/regTable[1][165] ), 
        .I2(\vrf/regTable[2][165] ), .I3(\vrf/regTable[3][165] ), .S0(n4780), 
        .S1(n4850), .ZN(n4066) );
  MUX4ND0BWP U6067 ( .I0(\vrf/regTable[4][165] ), .I1(\vrf/regTable[5][165] ), 
        .I2(\vrf/regTable[6][165] ), .I3(\vrf/regTable[7][165] ), .S0(n4780), 
        .S1(n4850), .ZN(n4067) );
  MUX2ND0BWP U6068 ( .I0(n4068), .I1(n4069), .S(n4901), .ZN(vectorData1[98])
         );
  MUX4ND0BWP U6069 ( .I0(\vrf/regTable[0][98] ), .I1(\vrf/regTable[1][98] ), 
        .I2(\vrf/regTable[2][98] ), .I3(\vrf/regTable[3][98] ), .S0(n4769), 
        .S1(n4839), .ZN(n4068) );
  MUX4ND0BWP U6070 ( .I0(\vrf/regTable[4][98] ), .I1(\vrf/regTable[5][98] ), 
        .I2(\vrf/regTable[6][98] ), .I3(\vrf/regTable[7][98] ), .S0(n4769), 
        .S1(n4839), .ZN(n4069) );
  MUX2ND0BWP U6071 ( .I0(n4070), .I1(n4071), .S(n4895), .ZN(vectorData1[34])
         );
  MUX4ND0BWP U6072 ( .I0(\vrf/regTable[0][34] ), .I1(\vrf/regTable[1][34] ), 
        .I2(\vrf/regTable[2][34] ), .I3(\vrf/regTable[3][34] ), .S0(n4758), 
        .S1(n4828), .ZN(n4070) );
  MUX4ND0BWP U6073 ( .I0(\vrf/regTable[4][34] ), .I1(\vrf/regTable[5][34] ), 
        .I2(\vrf/regTable[6][34] ), .I3(\vrf/regTable[7][34] ), .S0(n4758), 
        .S1(n4828), .ZN(n4071) );
  MUX2ND0BWP U6074 ( .I0(n4072), .I1(n4073), .S(n4906), .ZN(vectorData1[162])
         );
  MUX4ND0BWP U6075 ( .I0(\vrf/regTable[0][162] ), .I1(\vrf/regTable[1][162] ), 
        .I2(\vrf/regTable[2][162] ), .I3(\vrf/regTable[3][162] ), .S0(n4780), 
        .S1(n4850), .ZN(n4072) );
  MUX4ND0BWP U6076 ( .I0(\vrf/regTable[4][162] ), .I1(\vrf/regTable[5][162] ), 
        .I2(\vrf/regTable[6][162] ), .I3(\vrf/regTable[7][162] ), .S0(n4780), 
        .S1(n4850), .ZN(n4073) );
  MUX2ND0BWP U6077 ( .I0(n4074), .I1(n4075), .S(n4901), .ZN(vectorData1[99])
         );
  MUX4ND0BWP U6078 ( .I0(\vrf/regTable[0][99] ), .I1(\vrf/regTable[1][99] ), 
        .I2(\vrf/regTable[2][99] ), .I3(\vrf/regTable[3][99] ), .S0(n4769), 
        .S1(n4839), .ZN(n4074) );
  MUX4ND0BWP U6079 ( .I0(\vrf/regTable[4][99] ), .I1(\vrf/regTable[5][99] ), 
        .I2(\vrf/regTable[6][99] ), .I3(\vrf/regTable[7][99] ), .S0(n4769), 
        .S1(n4839), .ZN(n4075) );
  MUX2ND0BWP U6080 ( .I0(n4076), .I1(n4077), .S(n4895), .ZN(vectorData1[35])
         );
  MUX4ND0BWP U6081 ( .I0(\vrf/regTable[0][35] ), .I1(\vrf/regTable[1][35] ), 
        .I2(\vrf/regTable[2][35] ), .I3(\vrf/regTable[3][35] ), .S0(n4758), 
        .S1(n4828), .ZN(n4076) );
  MUX4ND0BWP U6082 ( .I0(\vrf/regTable[4][35] ), .I1(\vrf/regTable[5][35] ), 
        .I2(\vrf/regTable[6][35] ), .I3(\vrf/regTable[7][35] ), .S0(n4758), 
        .S1(n4828), .ZN(n4077) );
  MUX2ND0BWP U6083 ( .I0(n4078), .I1(n4079), .S(n4906), .ZN(vectorData1[163])
         );
  MUX4ND0BWP U6084 ( .I0(\vrf/regTable[0][163] ), .I1(\vrf/regTable[1][163] ), 
        .I2(\vrf/regTable[2][163] ), .I3(\vrf/regTable[3][163] ), .S0(n4780), 
        .S1(n4850), .ZN(n4078) );
  MUX4ND0BWP U6085 ( .I0(\vrf/regTable[4][163] ), .I1(\vrf/regTable[5][163] ), 
        .I2(\vrf/regTable[6][163] ), .I3(\vrf/regTable[7][163] ), .S0(n4780), 
        .S1(n4850), .ZN(n4079) );
  MUX2ND0BWP U6086 ( .I0(n4080), .I1(n4081), .S(n4901), .ZN(vectorData1[100])
         );
  MUX4ND0BWP U6087 ( .I0(\vrf/regTable[0][100] ), .I1(\vrf/regTable[1][100] ), 
        .I2(\vrf/regTable[2][100] ), .I3(\vrf/regTable[3][100] ), .S0(n4769), 
        .S1(n4839), .ZN(n4080) );
  MUX4ND0BWP U6088 ( .I0(\vrf/regTable[4][100] ), .I1(\vrf/regTable[5][100] ), 
        .I2(\vrf/regTable[6][100] ), .I3(\vrf/regTable[7][100] ), .S0(n4769), 
        .S1(n4839), .ZN(n4081) );
  MUX2ND0BWP U6089 ( .I0(n4082), .I1(n4083), .S(n4896), .ZN(vectorData1[36])
         );
  MUX4ND0BWP U6090 ( .I0(\vrf/regTable[0][36] ), .I1(\vrf/regTable[1][36] ), 
        .I2(\vrf/regTable[2][36] ), .I3(\vrf/regTable[3][36] ), .S0(n4759), 
        .S1(n4829), .ZN(n4082) );
  MUX4ND0BWP U6091 ( .I0(\vrf/regTable[4][36] ), .I1(\vrf/regTable[5][36] ), 
        .I2(\vrf/regTable[6][36] ), .I3(\vrf/regTable[7][36] ), .S0(n4759), 
        .S1(n4829), .ZN(n4083) );
  MUX2ND0BWP U6092 ( .I0(n4084), .I1(n4085), .S(n4906), .ZN(vectorData1[164])
         );
  MUX4ND0BWP U6093 ( .I0(\vrf/regTable[0][164] ), .I1(\vrf/regTable[1][164] ), 
        .I2(\vrf/regTable[2][164] ), .I3(\vrf/regTable[3][164] ), .S0(n4780), 
        .S1(n4850), .ZN(n4084) );
  MUX4ND0BWP U6094 ( .I0(\vrf/regTable[4][164] ), .I1(\vrf/regTable[5][164] ), 
        .I2(\vrf/regTable[6][164] ), .I3(\vrf/regTable[7][164] ), .S0(n4780), 
        .S1(n4850), .ZN(n4085) );
  MUX2ND0BWP U6095 ( .I0(n4086), .I1(n4087), .S(n5082), .ZN(vectorData2[179])
         );
  MUX4ND0BWP U6096 ( .I0(\vrf/regTable[0][179] ), .I1(\vrf/regTable[1][179] ), 
        .I2(\vrf/regTable[2][179] ), .I3(\vrf/regTable[3][179] ), .S0(n4957), 
        .S1(n5027), .ZN(n4086) );
  MUX4ND0BWP U6097 ( .I0(\vrf/regTable[4][179] ), .I1(\vrf/regTable[5][179] ), 
        .I2(\vrf/regTable[6][179] ), .I3(\vrf/regTable[7][179] ), .S0(n4957), 
        .S1(n5027), .ZN(n4087) );
  MUX2ND0BWP U6098 ( .I0(n4088), .I1(n4089), .S(n5083), .ZN(vectorData2[180])
         );
  MUX4ND0BWP U6099 ( .I0(\vrf/regTable[0][180] ), .I1(\vrf/regTable[1][180] ), 
        .I2(\vrf/regTable[2][180] ), .I3(\vrf/regTable[3][180] ), .S0(n4958), 
        .S1(n5028), .ZN(n4088) );
  MUX4ND0BWP U6100 ( .I0(\vrf/regTable[4][180] ), .I1(\vrf/regTable[5][180] ), 
        .I2(\vrf/regTable[6][180] ), .I3(\vrf/regTable[7][180] ), .S0(n4958), 
        .S1(n5028), .ZN(n4089) );
  MUX2ND0BWP U6101 ( .I0(n4090), .I1(n4091), .S(n5078), .ZN(vectorData2[128])
         );
  MUX4ND0BWP U6102 ( .I0(\vrf/regTable[0][128] ), .I1(\vrf/regTable[1][128] ), 
        .I2(\vrf/regTable[2][128] ), .I3(\vrf/regTable[3][128] ), .S0(n4949), 
        .S1(n5019), .ZN(n4090) );
  MUX4ND0BWP U6103 ( .I0(\vrf/regTable[4][128] ), .I1(\vrf/regTable[5][128] ), 
        .I2(\vrf/regTable[6][128] ), .I3(\vrf/regTable[7][128] ), .S0(n4949), 
        .S1(n5019), .ZN(n4091) );
  MUX2ND0BWP U6104 ( .I0(n4092), .I1(n4093), .S(n5078), .ZN(vectorData2[129])
         );
  MUX4ND0BWP U6105 ( .I0(\vrf/regTable[0][129] ), .I1(\vrf/regTable[1][129] ), 
        .I2(\vrf/regTable[2][129] ), .I3(\vrf/regTable[3][129] ), .S0(n4949), 
        .S1(n5019), .ZN(n4092) );
  MUX4ND0BWP U6106 ( .I0(\vrf/regTable[4][129] ), .I1(\vrf/regTable[5][129] ), 
        .I2(\vrf/regTable[6][129] ), .I3(\vrf/regTable[7][129] ), .S0(n4949), 
        .S1(n5019), .ZN(n4093) );
  MUX2ND0BWP U6107 ( .I0(n4094), .I1(n4095), .S(n5078), .ZN(vectorData2[130])
         );
  MUX4ND0BWP U6108 ( .I0(\vrf/regTable[0][130] ), .I1(\vrf/regTable[1][130] ), 
        .I2(\vrf/regTable[2][130] ), .I3(\vrf/regTable[3][130] ), .S0(n4949), 
        .S1(n5019), .ZN(n4094) );
  MUX4ND0BWP U6109 ( .I0(\vrf/regTable[4][130] ), .I1(\vrf/regTable[5][130] ), 
        .I2(\vrf/regTable[6][130] ), .I3(\vrf/regTable[7][130] ), .S0(n4949), 
        .S1(n5019), .ZN(n4095) );
  MUX2ND0BWP U6110 ( .I0(n4096), .I1(n4097), .S(n5079), .ZN(vectorData2[133])
         );
  MUX4ND0BWP U6111 ( .I0(\vrf/regTable[0][133] ), .I1(\vrf/regTable[1][133] ), 
        .I2(\vrf/regTable[2][133] ), .I3(\vrf/regTable[3][133] ), .S0(n4950), 
        .S1(n5020), .ZN(n4096) );
  MUX4ND0BWP U6112 ( .I0(\vrf/regTable[4][133] ), .I1(\vrf/regTable[5][133] ), 
        .I2(\vrf/regTable[6][133] ), .I3(\vrf/regTable[7][133] ), .S0(n4950), 
        .S1(n5020), .ZN(n4097) );
  MUX2ND0BWP U6113 ( .I0(n4098), .I1(n4099), .S(n5079), .ZN(vectorData2[134])
         );
  MUX4ND0BWP U6114 ( .I0(\vrf/regTable[0][134] ), .I1(\vrf/regTable[1][134] ), 
        .I2(\vrf/regTable[2][134] ), .I3(\vrf/regTable[3][134] ), .S0(n4950), 
        .S1(n5020), .ZN(n4098) );
  MUX4ND0BWP U6115 ( .I0(\vrf/regTable[4][134] ), .I1(\vrf/regTable[5][134] ), 
        .I2(\vrf/regTable[6][134] ), .I3(\vrf/regTable[7][134] ), .S0(n4950), 
        .S1(n5020), .ZN(n4099) );
  MUX2ND0BWP U6116 ( .I0(n4100), .I1(n4101), .S(n5079), .ZN(vectorData2[135])
         );
  MUX4ND0BWP U6117 ( .I0(\vrf/regTable[0][135] ), .I1(\vrf/regTable[1][135] ), 
        .I2(\vrf/regTable[2][135] ), .I3(\vrf/regTable[3][135] ), .S0(n4950), 
        .S1(n5020), .ZN(n4100) );
  MUX4ND0BWP U6118 ( .I0(\vrf/regTable[4][135] ), .I1(\vrf/regTable[5][135] ), 
        .I2(\vrf/regTable[6][135] ), .I3(\vrf/regTable[7][135] ), .S0(n4950), 
        .S1(n5020), .ZN(n4101) );
  MUX2ND0BWP U6119 ( .I0(n4102), .I1(n4103), .S(n5079), .ZN(vectorData2[136])
         );
  MUX4ND0BWP U6120 ( .I0(\vrf/regTable[0][136] ), .I1(\vrf/regTable[1][136] ), 
        .I2(\vrf/regTable[2][136] ), .I3(\vrf/regTable[3][136] ), .S0(n4950), 
        .S1(n5020), .ZN(n4102) );
  MUX4ND0BWP U6121 ( .I0(\vrf/regTable[4][136] ), .I1(\vrf/regTable[5][136] ), 
        .I2(\vrf/regTable[6][136] ), .I3(\vrf/regTable[7][136] ), .S0(n4950), 
        .S1(n5020), .ZN(n4103) );
  MUX2ND0BWP U6122 ( .I0(n4104), .I1(n4105), .S(n5079), .ZN(vectorData2[137])
         );
  MUX4ND0BWP U6123 ( .I0(\vrf/regTable[0][137] ), .I1(\vrf/regTable[1][137] ), 
        .I2(\vrf/regTable[2][137] ), .I3(\vrf/regTable[3][137] ), .S0(n4950), 
        .S1(n5020), .ZN(n4104) );
  MUX4ND0BWP U6124 ( .I0(\vrf/regTable[4][137] ), .I1(\vrf/regTable[5][137] ), 
        .I2(\vrf/regTable[6][137] ), .I3(\vrf/regTable[7][137] ), .S0(n4950), 
        .S1(n5020), .ZN(n4105) );
  MUX2ND0BWP U6125 ( .I0(n4106), .I1(n4107), .S(n5079), .ZN(vectorData2[138])
         );
  MUX4ND0BWP U6126 ( .I0(\vrf/regTable[0][138] ), .I1(\vrf/regTable[1][138] ), 
        .I2(\vrf/regTable[2][138] ), .I3(\vrf/regTable[3][138] ), .S0(n4951), 
        .S1(n5021), .ZN(n4106) );
  MUX4ND0BWP U6127 ( .I0(\vrf/regTable[4][138] ), .I1(\vrf/regTable[5][138] ), 
        .I2(\vrf/regTable[6][138] ), .I3(\vrf/regTable[7][138] ), .S0(n4951), 
        .S1(n5021), .ZN(n4107) );
  MUX2ND0BWP U6128 ( .I0(n4108), .I1(n4109), .S(n5079), .ZN(vectorData2[139])
         );
  MUX4ND0BWP U6129 ( .I0(\vrf/regTable[0][139] ), .I1(\vrf/regTable[1][139] ), 
        .I2(\vrf/regTable[2][139] ), .I3(\vrf/regTable[3][139] ), .S0(n4951), 
        .S1(n5021), .ZN(n4108) );
  MUX4ND0BWP U6130 ( .I0(\vrf/regTable[4][139] ), .I1(\vrf/regTable[5][139] ), 
        .I2(\vrf/regTable[6][139] ), .I3(\vrf/regTable[7][139] ), .S0(n4951), 
        .S1(n5021), .ZN(n4109) );
  MUX2ND0BWP U6131 ( .I0(n4110), .I1(n4111), .S(n5079), .ZN(vectorData2[140])
         );
  MUX4ND0BWP U6132 ( .I0(\vrf/regTable[0][140] ), .I1(\vrf/regTable[1][140] ), 
        .I2(\vrf/regTable[2][140] ), .I3(\vrf/regTable[3][140] ), .S0(n4951), 
        .S1(n5021), .ZN(n4110) );
  MUX4ND0BWP U6133 ( .I0(\vrf/regTable[4][140] ), .I1(\vrf/regTable[5][140] ), 
        .I2(\vrf/regTable[6][140] ), .I3(\vrf/regTable[7][140] ), .S0(n4951), 
        .S1(n5021), .ZN(n4111) );
  MUX2ND0BWP U6134 ( .I0(n4112), .I1(n4113), .S(n5079), .ZN(vectorData2[141])
         );
  MUX4ND0BWP U6135 ( .I0(\vrf/regTable[0][141] ), .I1(\vrf/regTable[1][141] ), 
        .I2(\vrf/regTable[2][141] ), .I3(\vrf/regTable[3][141] ), .S0(n4951), 
        .S1(n5021), .ZN(n4112) );
  MUX4ND0BWP U6136 ( .I0(\vrf/regTable[4][141] ), .I1(\vrf/regTable[5][141] ), 
        .I2(\vrf/regTable[6][141] ), .I3(\vrf/regTable[7][141] ), .S0(n4951), 
        .S1(n5021), .ZN(n4113) );
  MUX2ND0BWP U6137 ( .I0(n4114), .I1(n4115), .S(n5079), .ZN(vectorData2[142])
         );
  MUX4ND0BWP U6138 ( .I0(\vrf/regTable[0][142] ), .I1(\vrf/regTable[1][142] ), 
        .I2(\vrf/regTable[2][142] ), .I3(\vrf/regTable[3][142] ), .S0(n4951), 
        .S1(n5021), .ZN(n4114) );
  MUX4ND0BWP U6139 ( .I0(\vrf/regTable[4][142] ), .I1(\vrf/regTable[5][142] ), 
        .I2(\vrf/regTable[6][142] ), .I3(\vrf/regTable[7][142] ), .S0(n4951), 
        .S1(n5021), .ZN(n4115) );
  MUX2ND0BWP U6140 ( .I0(n4116), .I1(n4117), .S(n5079), .ZN(vectorData2[143])
         );
  MUX4ND0BWP U6141 ( .I0(\vrf/regTable[0][143] ), .I1(\vrf/regTable[1][143] ), 
        .I2(\vrf/regTable[2][143] ), .I3(\vrf/regTable[3][143] ), .S0(n4951), 
        .S1(n5021), .ZN(n4116) );
  MUX4ND0BWP U6142 ( .I0(\vrf/regTable[4][143] ), .I1(\vrf/regTable[5][143] ), 
        .I2(\vrf/regTable[6][143] ), .I3(\vrf/regTable[7][143] ), .S0(n4951), 
        .S1(n5021), .ZN(n4117) );
  MUX2ND0BWP U6143 ( .I0(n4118), .I1(n4119), .S(n5088), .ZN(vectorData2[240])
         );
  MUX4ND0BWP U6144 ( .I0(\vrf/regTable[0][240] ), .I1(\vrf/regTable[1][240] ), 
        .I2(\vrf/regTable[2][240] ), .I3(\vrf/regTable[3][240] ), .S0(n4968), 
        .S1(n5038), .ZN(n4118) );
  MUX4ND0BWP U6145 ( .I0(\vrf/regTable[4][240] ), .I1(\vrf/regTable[5][240] ), 
        .I2(\vrf/regTable[6][240] ), .I3(\vrf/regTable[7][240] ), .S0(n4968), 
        .S1(n5038), .ZN(n4119) );
  MUX2ND0BWP U6146 ( .I0(n4120), .I1(n4121), .S(n5088), .ZN(vectorData2[241])
         );
  MUX4ND0BWP U6147 ( .I0(\vrf/regTable[0][241] ), .I1(\vrf/regTable[1][241] ), 
        .I2(\vrf/regTable[2][241] ), .I3(\vrf/regTable[3][241] ), .S0(n4968), 
        .S1(n5038), .ZN(n4120) );
  MUX4ND0BWP U6148 ( .I0(\vrf/regTable[4][241] ), .I1(\vrf/regTable[5][241] ), 
        .I2(\vrf/regTable[6][241] ), .I3(\vrf/regTable[7][241] ), .S0(n4968), 
        .S1(n5038), .ZN(n4121) );
  MUX2ND0BWP U6149 ( .I0(n4122), .I1(n4123), .S(n5088), .ZN(vectorData2[242])
         );
  MUX4ND0BWP U6150 ( .I0(\vrf/regTable[0][242] ), .I1(\vrf/regTable[1][242] ), 
        .I2(\vrf/regTable[2][242] ), .I3(\vrf/regTable[3][242] ), .S0(n4968), 
        .S1(n5038), .ZN(n4122) );
  MUX4ND0BWP U6151 ( .I0(\vrf/regTable[4][242] ), .I1(\vrf/regTable[5][242] ), 
        .I2(\vrf/regTable[6][242] ), .I3(\vrf/regTable[7][242] ), .S0(n4968), 
        .S1(n5038), .ZN(n4123) );
  MUX2ND0BWP U6152 ( .I0(n4124), .I1(n4125), .S(n5088), .ZN(vectorData2[245])
         );
  MUX4ND0BWP U6153 ( .I0(\vrf/regTable[0][245] ), .I1(\vrf/regTable[1][245] ), 
        .I2(\vrf/regTable[2][245] ), .I3(\vrf/regTable[3][245] ), .S0(n4968), 
        .S1(n5038), .ZN(n4124) );
  MUX4ND0BWP U6154 ( .I0(\vrf/regTable[4][245] ), .I1(\vrf/regTable[5][245] ), 
        .I2(\vrf/regTable[6][245] ), .I3(\vrf/regTable[7][245] ), .S0(n4968), 
        .S1(n5038), .ZN(n4125) );
  MUX2ND0BWP U6155 ( .I0(n4126), .I1(n4127), .S(n5088), .ZN(vectorData2[246])
         );
  MUX4ND0BWP U6156 ( .I0(\vrf/regTable[0][246] ), .I1(\vrf/regTable[1][246] ), 
        .I2(\vrf/regTable[2][246] ), .I3(\vrf/regTable[3][246] ), .S0(n4969), 
        .S1(n5039), .ZN(n4126) );
  MUX4ND0BWP U6157 ( .I0(\vrf/regTable[4][246] ), .I1(\vrf/regTable[5][246] ), 
        .I2(\vrf/regTable[6][246] ), .I3(\vrf/regTable[7][246] ), .S0(n4969), 
        .S1(n5039), .ZN(n4127) );
  MUX2ND0BWP U6158 ( .I0(n4128), .I1(n4129), .S(n5088), .ZN(vectorData2[247])
         );
  MUX4ND0BWP U6159 ( .I0(\vrf/regTable[0][247] ), .I1(\vrf/regTable[1][247] ), 
        .I2(\vrf/regTable[2][247] ), .I3(\vrf/regTable[3][247] ), .S0(n4969), 
        .S1(n5039), .ZN(n4128) );
  MUX4ND0BWP U6160 ( .I0(\vrf/regTable[4][247] ), .I1(\vrf/regTable[5][247] ), 
        .I2(\vrf/regTable[6][247] ), .I3(\vrf/regTable[7][247] ), .S0(n4969), 
        .S1(n5039), .ZN(n4129) );
  MUX2ND0BWP U6161 ( .I0(n4130), .I1(n4131), .S(n5088), .ZN(vectorData2[248])
         );
  MUX4ND0BWP U6162 ( .I0(\vrf/regTable[0][248] ), .I1(\vrf/regTable[1][248] ), 
        .I2(\vrf/regTable[2][248] ), .I3(\vrf/regTable[3][248] ), .S0(n4969), 
        .S1(n5039), .ZN(n4130) );
  MUX4ND0BWP U6163 ( .I0(\vrf/regTable[4][248] ), .I1(\vrf/regTable[5][248] ), 
        .I2(\vrf/regTable[6][248] ), .I3(\vrf/regTable[7][248] ), .S0(n4969), 
        .S1(n5039), .ZN(n4131) );
  MUX2ND0BWP U6164 ( .I0(n4132), .I1(n4133), .S(n5088), .ZN(vectorData2[249])
         );
  MUX4ND0BWP U6165 ( .I0(\vrf/regTable[0][249] ), .I1(\vrf/regTable[1][249] ), 
        .I2(\vrf/regTable[2][249] ), .I3(\vrf/regTable[3][249] ), .S0(n4969), 
        .S1(n5039), .ZN(n4132) );
  MUX4ND0BWP U6166 ( .I0(\vrf/regTable[4][249] ), .I1(\vrf/regTable[5][249] ), 
        .I2(\vrf/regTable[6][249] ), .I3(\vrf/regTable[7][249] ), .S0(n4969), 
        .S1(n5039), .ZN(n4133) );
  MUX2ND0BWP U6167 ( .I0(n4134), .I1(n4135), .S(n5088), .ZN(vectorData2[250])
         );
  MUX4ND0BWP U6168 ( .I0(\vrf/regTable[0][250] ), .I1(\vrf/regTable[1][250] ), 
        .I2(\vrf/regTable[2][250] ), .I3(\vrf/regTable[3][250] ), .S0(n4969), 
        .S1(n5039), .ZN(n4134) );
  MUX4ND0BWP U6169 ( .I0(\vrf/regTable[4][250] ), .I1(\vrf/regTable[5][250] ), 
        .I2(\vrf/regTable[6][250] ), .I3(\vrf/regTable[7][250] ), .S0(n4969), 
        .S1(n5039), .ZN(n4135) );
  MUX2ND0BWP U6170 ( .I0(n4136), .I1(n4137), .S(n5088), .ZN(vectorData2[251])
         );
  MUX4ND0BWP U6171 ( .I0(\vrf/regTable[0][251] ), .I1(\vrf/regTable[1][251] ), 
        .I2(\vrf/regTable[2][251] ), .I3(\vrf/regTable[3][251] ), .S0(n4969), 
        .S1(n5039), .ZN(n4136) );
  MUX4ND0BWP U6172 ( .I0(\vrf/regTable[4][251] ), .I1(\vrf/regTable[5][251] ), 
        .I2(\vrf/regTable[6][251] ), .I3(\vrf/regTable[7][251] ), .S0(n4969), 
        .S1(n5039), .ZN(n4137) );
  MUX2ND0BWP U6173 ( .I0(n4138), .I1(n4139), .S(n5089), .ZN(vectorData2[252])
         );
  MUX4ND0BWP U6174 ( .I0(\vrf/regTable[0][252] ), .I1(\vrf/regTable[1][252] ), 
        .I2(\vrf/regTable[2][252] ), .I3(\vrf/regTable[3][252] ), .S0(n4970), 
        .S1(n5040), .ZN(n4138) );
  MUX4ND0BWP U6175 ( .I0(\vrf/regTable[4][252] ), .I1(\vrf/regTable[5][252] ), 
        .I2(\vrf/regTable[6][252] ), .I3(\vrf/regTable[7][252] ), .S0(n4970), 
        .S1(n5040), .ZN(n4139) );
  MUX2ND0BWP U6176 ( .I0(n4140), .I1(n4141), .S(n5089), .ZN(vectorData2[253])
         );
  MUX4ND0BWP U6177 ( .I0(\vrf/regTable[0][253] ), .I1(\vrf/regTable[1][253] ), 
        .I2(\vrf/regTable[2][253] ), .I3(\vrf/regTable[3][253] ), .S0(n4970), 
        .S1(n5040), .ZN(n4140) );
  MUX4ND0BWP U6178 ( .I0(\vrf/regTable[4][253] ), .I1(\vrf/regTable[5][253] ), 
        .I2(\vrf/regTable[6][253] ), .I3(\vrf/regTable[7][253] ), .S0(n4970), 
        .S1(n5040), .ZN(n4141) );
  MUX2ND0BWP U6179 ( .I0(n4142), .I1(n4143), .S(n5089), .ZN(vectorData2[254])
         );
  MUX4ND0BWP U6180 ( .I0(\vrf/regTable[0][254] ), .I1(\vrf/regTable[1][254] ), 
        .I2(\vrf/regTable[2][254] ), .I3(\vrf/regTable[3][254] ), .S0(n4970), 
        .S1(n5040), .ZN(n4142) );
  MUX4ND0BWP U6181 ( .I0(\vrf/regTable[4][254] ), .I1(\vrf/regTable[5][254] ), 
        .I2(\vrf/regTable[6][254] ), .I3(\vrf/regTable[7][254] ), .S0(n4970), 
        .S1(n5040), .ZN(n4143) );
  MUX2ND0BWP U6182 ( .I0(n4144), .I1(n4145), .S(n5089), .ZN(vectorData2[255])
         );
  MUX4ND0BWP U6183 ( .I0(\vrf/regTable[0][255] ), .I1(\vrf/regTable[1][255] ), 
        .I2(\vrf/regTable[2][255] ), .I3(\vrf/regTable[3][255] ), .S0(n4970), 
        .S1(n5040), .ZN(n4144) );
  MUX4ND0BWP U6184 ( .I0(\vrf/regTable[4][255] ), .I1(\vrf/regTable[5][255] ), 
        .I2(\vrf/regTable[6][255] ), .I3(\vrf/regTable[7][255] ), .S0(n4970), 
        .S1(n5040), .ZN(n4145) );
  MUX2ND0BWP U6185 ( .I0(n4146), .I1(n4147), .S(n5078), .ZN(vectorData2[131])
         );
  MUX4ND0BWP U6186 ( .I0(\vrf/regTable[0][131] ), .I1(\vrf/regTable[1][131] ), 
        .I2(\vrf/regTable[2][131] ), .I3(\vrf/regTable[3][131] ), .S0(n4949), 
        .S1(n5019), .ZN(n4146) );
  MUX4ND0BWP U6187 ( .I0(\vrf/regTable[4][131] ), .I1(\vrf/regTable[5][131] ), 
        .I2(\vrf/regTable[6][131] ), .I3(\vrf/regTable[7][131] ), .S0(n4949), 
        .S1(n5019), .ZN(n4147) );
  MUX2ND0BWP U6188 ( .I0(n4148), .I1(n4149), .S(n5088), .ZN(vectorData2[243])
         );
  MUX4ND0BWP U6189 ( .I0(\vrf/regTable[0][243] ), .I1(\vrf/regTable[1][243] ), 
        .I2(\vrf/regTable[2][243] ), .I3(\vrf/regTable[3][243] ), .S0(n4968), 
        .S1(n5038), .ZN(n4148) );
  MUX4ND0BWP U6190 ( .I0(\vrf/regTable[4][243] ), .I1(\vrf/regTable[5][243] ), 
        .I2(\vrf/regTable[6][243] ), .I3(\vrf/regTable[7][243] ), .S0(n4968), 
        .S1(n5038), .ZN(n4149) );
  MUX2ND0BWP U6191 ( .I0(n4150), .I1(n4151), .S(n5079), .ZN(vectorData2[132])
         );
  MUX4ND0BWP U6192 ( .I0(\vrf/regTable[0][132] ), .I1(\vrf/regTable[1][132] ), 
        .I2(\vrf/regTable[2][132] ), .I3(\vrf/regTable[3][132] ), .S0(n4950), 
        .S1(n5020), .ZN(n4150) );
  MUX4ND0BWP U6193 ( .I0(\vrf/regTable[4][132] ), .I1(\vrf/regTable[5][132] ), 
        .I2(\vrf/regTable[6][132] ), .I3(\vrf/regTable[7][132] ), .S0(n4950), 
        .S1(n5020), .ZN(n4151) );
  MUX2ND0BWP U6194 ( .I0(n4152), .I1(n4153), .S(n5088), .ZN(vectorData2[244])
         );
  MUX4ND0BWP U6195 ( .I0(\vrf/regTable[0][244] ), .I1(\vrf/regTable[1][244] ), 
        .I2(\vrf/regTable[2][244] ), .I3(\vrf/regTable[3][244] ), .S0(n4968), 
        .S1(n5038), .ZN(n4152) );
  MUX4ND0BWP U6196 ( .I0(\vrf/regTable[4][244] ), .I1(\vrf/regTable[5][244] ), 
        .I2(\vrf/regTable[6][244] ), .I3(\vrf/regTable[7][244] ), .S0(n4968), 
        .S1(n5038), .ZN(n4153) );
  MUX2ND0BWP U6197 ( .I0(n4154), .I1(n4155), .S(n5086), .ZN(vectorData2[224])
         );
  MUX4ND0BWP U6198 ( .I0(\vrf/regTable[0][224] ), .I1(\vrf/regTable[1][224] ), 
        .I2(\vrf/regTable[2][224] ), .I3(\vrf/regTable[3][224] ), .S0(n4965), 
        .S1(n5035), .ZN(n4154) );
  MUX4ND0BWP U6199 ( .I0(\vrf/regTable[4][224] ), .I1(\vrf/regTable[5][224] ), 
        .I2(\vrf/regTable[6][224] ), .I3(\vrf/regTable[7][224] ), .S0(n4965), 
        .S1(n5035), .ZN(n4155) );
  MUX2ND0BWP U6200 ( .I0(n4156), .I1(n4157), .S(n5086), .ZN(vectorData2[225])
         );
  MUX4ND0BWP U6201 ( .I0(\vrf/regTable[0][225] ), .I1(\vrf/regTable[1][225] ), 
        .I2(\vrf/regTable[2][225] ), .I3(\vrf/regTable[3][225] ), .S0(n4965), 
        .S1(n5035), .ZN(n4156) );
  MUX4ND0BWP U6202 ( .I0(\vrf/regTable[4][225] ), .I1(\vrf/regTable[5][225] ), 
        .I2(\vrf/regTable[6][225] ), .I3(\vrf/regTable[7][225] ), .S0(n4965), 
        .S1(n5035), .ZN(n4157) );
  MUX2ND0BWP U6203 ( .I0(n4158), .I1(n4159), .S(n5086), .ZN(vectorData2[226])
         );
  MUX4ND0BWP U6204 ( .I0(\vrf/regTable[0][226] ), .I1(\vrf/regTable[1][226] ), 
        .I2(\vrf/regTable[2][226] ), .I3(\vrf/regTable[3][226] ), .S0(n4965), 
        .S1(n5035), .ZN(n4158) );
  MUX4ND0BWP U6205 ( .I0(\vrf/regTable[4][226] ), .I1(\vrf/regTable[5][226] ), 
        .I2(\vrf/regTable[6][226] ), .I3(\vrf/regTable[7][226] ), .S0(n4965), 
        .S1(n5035), .ZN(n4159) );
  MUX2ND0BWP U6206 ( .I0(n4160), .I1(n4161), .S(n5087), .ZN(vectorData2[229])
         );
  MUX4ND0BWP U6207 ( .I0(\vrf/regTable[0][229] ), .I1(\vrf/regTable[1][229] ), 
        .I2(\vrf/regTable[2][229] ), .I3(\vrf/regTable[3][229] ), .S0(n4966), 
        .S1(n5036), .ZN(n4160) );
  MUX4ND0BWP U6208 ( .I0(\vrf/regTable[4][229] ), .I1(\vrf/regTable[5][229] ), 
        .I2(\vrf/regTable[6][229] ), .I3(\vrf/regTable[7][229] ), .S0(n4966), 
        .S1(n5036), .ZN(n4161) );
  MUX2ND0BWP U6209 ( .I0(n4162), .I1(n4163), .S(n5087), .ZN(vectorData2[230])
         );
  MUX4ND0BWP U6210 ( .I0(\vrf/regTable[0][230] ), .I1(\vrf/regTable[1][230] ), 
        .I2(\vrf/regTable[2][230] ), .I3(\vrf/regTable[3][230] ), .S0(n4966), 
        .S1(n5036), .ZN(n4162) );
  MUX4ND0BWP U6211 ( .I0(\vrf/regTable[4][230] ), .I1(\vrf/regTable[5][230] ), 
        .I2(\vrf/regTable[6][230] ), .I3(\vrf/regTable[7][230] ), .S0(n4966), 
        .S1(n5036), .ZN(n4163) );
  MUX2ND0BWP U6212 ( .I0(n4164), .I1(n4165), .S(n5087), .ZN(vectorData2[231])
         );
  MUX4ND0BWP U6213 ( .I0(\vrf/regTable[0][231] ), .I1(\vrf/regTable[1][231] ), 
        .I2(\vrf/regTable[2][231] ), .I3(\vrf/regTable[3][231] ), .S0(n4966), 
        .S1(n5036), .ZN(n4164) );
  MUX4ND0BWP U6214 ( .I0(\vrf/regTable[4][231] ), .I1(\vrf/regTable[5][231] ), 
        .I2(\vrf/regTable[6][231] ), .I3(\vrf/regTable[7][231] ), .S0(n4966), 
        .S1(n5036), .ZN(n4165) );
  MUX2ND0BWP U6215 ( .I0(n4166), .I1(n4167), .S(n5087), .ZN(vectorData2[232])
         );
  MUX4ND0BWP U6216 ( .I0(\vrf/regTable[0][232] ), .I1(\vrf/regTable[1][232] ), 
        .I2(\vrf/regTable[2][232] ), .I3(\vrf/regTable[3][232] ), .S0(n4966), 
        .S1(n5036), .ZN(n4166) );
  MUX4ND0BWP U6217 ( .I0(\vrf/regTable[4][232] ), .I1(\vrf/regTable[5][232] ), 
        .I2(\vrf/regTable[6][232] ), .I3(\vrf/regTable[7][232] ), .S0(n4966), 
        .S1(n5036), .ZN(n4167) );
  MUX2ND0BWP U6218 ( .I0(n4168), .I1(n4169), .S(n5087), .ZN(vectorData2[233])
         );
  MUX4ND0BWP U6219 ( .I0(\vrf/regTable[0][233] ), .I1(\vrf/regTable[1][233] ), 
        .I2(\vrf/regTable[2][233] ), .I3(\vrf/regTable[3][233] ), .S0(n4966), 
        .S1(n5036), .ZN(n4168) );
  MUX4ND0BWP U6220 ( .I0(\vrf/regTable[4][233] ), .I1(\vrf/regTable[5][233] ), 
        .I2(\vrf/regTable[6][233] ), .I3(\vrf/regTable[7][233] ), .S0(n4966), 
        .S1(n5036), .ZN(n4169) );
  MUX2ND0BWP U6221 ( .I0(n4170), .I1(n4171), .S(n5087), .ZN(vectorData2[234])
         );
  MUX4ND0BWP U6222 ( .I0(\vrf/regTable[0][234] ), .I1(\vrf/regTable[1][234] ), 
        .I2(\vrf/regTable[2][234] ), .I3(\vrf/regTable[3][234] ), .S0(n4967), 
        .S1(n5037), .ZN(n4170) );
  MUX4ND0BWP U6223 ( .I0(\vrf/regTable[4][234] ), .I1(\vrf/regTable[5][234] ), 
        .I2(\vrf/regTable[6][234] ), .I3(\vrf/regTable[7][234] ), .S0(n4967), 
        .S1(n5037), .ZN(n4171) );
  MUX2ND0BWP U6224 ( .I0(n4172), .I1(n4173), .S(n5087), .ZN(vectorData2[235])
         );
  MUX4ND0BWP U6225 ( .I0(\vrf/regTable[0][235] ), .I1(\vrf/regTable[1][235] ), 
        .I2(\vrf/regTable[2][235] ), .I3(\vrf/regTable[3][235] ), .S0(n4967), 
        .S1(n5037), .ZN(n4172) );
  MUX4ND0BWP U6226 ( .I0(\vrf/regTable[4][235] ), .I1(\vrf/regTable[5][235] ), 
        .I2(\vrf/regTable[6][235] ), .I3(\vrf/regTable[7][235] ), .S0(n4967), 
        .S1(n5037), .ZN(n4173) );
  MUX2ND0BWP U6227 ( .I0(n4174), .I1(n4175), .S(n5087), .ZN(vectorData2[236])
         );
  MUX4ND0BWP U6228 ( .I0(\vrf/regTable[0][236] ), .I1(\vrf/regTable[1][236] ), 
        .I2(\vrf/regTable[2][236] ), .I3(\vrf/regTable[3][236] ), .S0(n4967), 
        .S1(n5037), .ZN(n4174) );
  MUX4ND0BWP U6229 ( .I0(\vrf/regTable[4][236] ), .I1(\vrf/regTable[5][236] ), 
        .I2(\vrf/regTable[6][236] ), .I3(\vrf/regTable[7][236] ), .S0(n4967), 
        .S1(n5037), .ZN(n4175) );
  MUX2ND0BWP U6230 ( .I0(n4176), .I1(n4177), .S(n5087), .ZN(vectorData2[237])
         );
  MUX4ND0BWP U6231 ( .I0(\vrf/regTable[0][237] ), .I1(\vrf/regTable[1][237] ), 
        .I2(\vrf/regTable[2][237] ), .I3(\vrf/regTable[3][237] ), .S0(n4967), 
        .S1(n5037), .ZN(n4176) );
  MUX4ND0BWP U6232 ( .I0(\vrf/regTable[4][237] ), .I1(\vrf/regTable[5][237] ), 
        .I2(\vrf/regTable[6][237] ), .I3(\vrf/regTable[7][237] ), .S0(n4967), 
        .S1(n5037), .ZN(n4177) );
  MUX2ND0BWP U6233 ( .I0(n4178), .I1(n4179), .S(n5087), .ZN(vectorData2[238])
         );
  MUX4ND0BWP U6234 ( .I0(\vrf/regTable[0][238] ), .I1(\vrf/regTable[1][238] ), 
        .I2(\vrf/regTable[2][238] ), .I3(\vrf/regTable[3][238] ), .S0(n4967), 
        .S1(n5037), .ZN(n4178) );
  MUX4ND0BWP U6235 ( .I0(\vrf/regTable[4][238] ), .I1(\vrf/regTable[5][238] ), 
        .I2(\vrf/regTable[6][238] ), .I3(\vrf/regTable[7][238] ), .S0(n4967), 
        .S1(n5037), .ZN(n4179) );
  MUX2ND0BWP U6236 ( .I0(n4180), .I1(n4181), .S(n5087), .ZN(vectorData2[239])
         );
  MUX4ND0BWP U6237 ( .I0(\vrf/regTable[0][239] ), .I1(\vrf/regTable[1][239] ), 
        .I2(\vrf/regTable[2][239] ), .I3(\vrf/regTable[3][239] ), .S0(n4967), 
        .S1(n5037), .ZN(n4180) );
  MUX4ND0BWP U6238 ( .I0(\vrf/regTable[4][239] ), .I1(\vrf/regTable[5][239] ), 
        .I2(\vrf/regTable[6][239] ), .I3(\vrf/regTable[7][239] ), .S0(n4967), 
        .S1(n5037), .ZN(n4181) );
  MUX2ND0BWP U6239 ( .I0(n4182), .I1(n4183), .S(n4899), .ZN(vectorData1[80])
         );
  MUX4ND0BWP U6240 ( .I0(\vrf/regTable[0][80] ), .I1(\vrf/regTable[1][80] ), 
        .I2(\vrf/regTable[2][80] ), .I3(\vrf/regTable[3][80] ), .S0(n4766), 
        .S1(n4836), .ZN(n4182) );
  MUX4ND0BWP U6241 ( .I0(\vrf/regTable[4][80] ), .I1(\vrf/regTable[5][80] ), 
        .I2(\vrf/regTable[6][80] ), .I3(\vrf/regTable[7][80] ), .S0(n4766), 
        .S1(n4836), .ZN(n4183) );
  MUX2ND0BWP U6242 ( .I0(n4184), .I1(n4185), .S(n4894), .ZN(vectorData1[16])
         );
  MUX4ND0BWP U6243 ( .I0(\vrf/regTable[0][16] ), .I1(\vrf/regTable[1][16] ), 
        .I2(\vrf/regTable[2][16] ), .I3(\vrf/regTable[3][16] ), .S0(n4755), 
        .S1(n4825), .ZN(n4184) );
  MUX4ND0BWP U6244 ( .I0(\vrf/regTable[4][16] ), .I1(\vrf/regTable[5][16] ), 
        .I2(\vrf/regTable[6][16] ), .I3(\vrf/regTable[7][16] ), .S0(n4755), 
        .S1(n4825), .ZN(n4185) );
  MUX2ND0BWP U6245 ( .I0(n4186), .I1(n4187), .S(n4905), .ZN(vectorData1[144])
         );
  MUX4ND0BWP U6246 ( .I0(\vrf/regTable[0][144] ), .I1(\vrf/regTable[1][144] ), 
        .I2(\vrf/regTable[2][144] ), .I3(\vrf/regTable[3][144] ), .S0(n4777), 
        .S1(n4847), .ZN(n4186) );
  MUX4ND0BWP U6247 ( .I0(\vrf/regTable[4][144] ), .I1(\vrf/regTable[5][144] ), 
        .I2(\vrf/regTable[6][144] ), .I3(\vrf/regTable[7][144] ), .S0(n4777), 
        .S1(n4847), .ZN(n4187) );
  MUX2ND0BWP U6248 ( .I0(n4188), .I1(n4189), .S(n4900), .ZN(vectorData1[95])
         );
  MUX4ND0BWP U6249 ( .I0(\vrf/regTable[0][95] ), .I1(\vrf/regTable[1][95] ), 
        .I2(\vrf/regTable[2][95] ), .I3(\vrf/regTable[3][95] ), .S0(n4768), 
        .S1(n4838), .ZN(n4188) );
  MUX4ND0BWP U6250 ( .I0(\vrf/regTable[4][95] ), .I1(\vrf/regTable[5][95] ), 
        .I2(\vrf/regTable[6][95] ), .I3(\vrf/regTable[7][95] ), .S0(n4768), 
        .S1(n4838), .ZN(n4189) );
  MUX2ND0BWP U6251 ( .I0(n4190), .I1(n4191), .S(n4895), .ZN(vectorData1[31])
         );
  MUX4ND0BWP U6252 ( .I0(\vrf/regTable[0][31] ), .I1(\vrf/regTable[1][31] ), 
        .I2(\vrf/regTable[2][31] ), .I3(\vrf/regTable[3][31] ), .S0(n4758), 
        .S1(n4828), .ZN(n4190) );
  MUX4ND0BWP U6253 ( .I0(\vrf/regTable[4][31] ), .I1(\vrf/regTable[5][31] ), 
        .I2(\vrf/regTable[6][31] ), .I3(\vrf/regTable[7][31] ), .S0(n4758), 
        .S1(n4828), .ZN(n4191) );
  MUX2ND0BWP U6254 ( .I0(n4192), .I1(n4193), .S(n4906), .ZN(vectorData1[159])
         );
  MUX4ND0BWP U6255 ( .I0(\vrf/regTable[0][159] ), .I1(\vrf/regTable[1][159] ), 
        .I2(\vrf/regTable[2][159] ), .I3(\vrf/regTable[3][159] ), .S0(n4779), 
        .S1(n4849), .ZN(n4192) );
  MUX4ND0BWP U6256 ( .I0(\vrf/regTable[4][159] ), .I1(\vrf/regTable[5][159] ), 
        .I2(\vrf/regTable[6][159] ), .I3(\vrf/regTable[7][159] ), .S0(n4779), 
        .S1(n4849), .ZN(n4193) );
  MUX2ND0BWP U6257 ( .I0(n4194), .I1(n4195), .S(n4900), .ZN(vectorData1[94])
         );
  MUX4ND0BWP U6258 ( .I0(\vrf/regTable[0][94] ), .I1(\vrf/regTable[1][94] ), 
        .I2(\vrf/regTable[2][94] ), .I3(\vrf/regTable[3][94] ), .S0(n4768), 
        .S1(n4838), .ZN(n4194) );
  MUX4ND0BWP U6259 ( .I0(\vrf/regTable[4][94] ), .I1(\vrf/regTable[5][94] ), 
        .I2(\vrf/regTable[6][94] ), .I3(\vrf/regTable[7][94] ), .S0(n4768), 
        .S1(n4838), .ZN(n4195) );
  MUX2ND0BWP U6260 ( .I0(n4196), .I1(n4197), .S(n4895), .ZN(vectorData1[30])
         );
  MUX4ND0BWP U6261 ( .I0(\vrf/regTable[0][30] ), .I1(\vrf/regTable[1][30] ), 
        .I2(\vrf/regTable[2][30] ), .I3(\vrf/regTable[3][30] ), .S0(n4758), 
        .S1(n4828), .ZN(n4196) );
  MUX4ND0BWP U6262 ( .I0(\vrf/regTable[4][30] ), .I1(\vrf/regTable[5][30] ), 
        .I2(\vrf/regTable[6][30] ), .I3(\vrf/regTable[7][30] ), .S0(n4758), 
        .S1(n4828), .ZN(n4197) );
  MUX2ND0BWP U6263 ( .I0(n4198), .I1(n4199), .S(n4906), .ZN(vectorData1[158])
         );
  MUX4ND0BWP U6264 ( .I0(\vrf/regTable[0][158] ), .I1(\vrf/regTable[1][158] ), 
        .I2(\vrf/regTable[2][158] ), .I3(\vrf/regTable[3][158] ), .S0(n4779), 
        .S1(n4849), .ZN(n4198) );
  MUX4ND0BWP U6265 ( .I0(\vrf/regTable[4][158] ), .I1(\vrf/regTable[5][158] ), 
        .I2(\vrf/regTable[6][158] ), .I3(\vrf/regTable[7][158] ), .S0(n4779), 
        .S1(n4849), .ZN(n4199) );
  MUX2ND0BWP U6266 ( .I0(n4200), .I1(n4201), .S(n4900), .ZN(vectorData1[93])
         );
  MUX4ND0BWP U6267 ( .I0(\vrf/regTable[0][93] ), .I1(\vrf/regTable[1][93] ), 
        .I2(\vrf/regTable[2][93] ), .I3(\vrf/regTable[3][93] ), .S0(n4768), 
        .S1(n4838), .ZN(n4200) );
  MUX4ND0BWP U6268 ( .I0(\vrf/regTable[4][93] ), .I1(\vrf/regTable[5][93] ), 
        .I2(\vrf/regTable[6][93] ), .I3(\vrf/regTable[7][93] ), .S0(n4768), 
        .S1(n4838), .ZN(n4201) );
  MUX2ND0BWP U6269 ( .I0(n4202), .I1(n4203), .S(n4895), .ZN(vectorData1[29])
         );
  MUX4ND0BWP U6270 ( .I0(\vrf/regTable[0][29] ), .I1(\vrf/regTable[1][29] ), 
        .I2(\vrf/regTable[2][29] ), .I3(\vrf/regTable[3][29] ), .S0(n4757), 
        .S1(n4827), .ZN(n4202) );
  MUX4ND0BWP U6271 ( .I0(\vrf/regTable[4][29] ), .I1(\vrf/regTable[5][29] ), 
        .I2(\vrf/regTable[6][29] ), .I3(\vrf/regTable[7][29] ), .S0(n4757), 
        .S1(n4827), .ZN(n4203) );
  MUX2ND0BWP U6272 ( .I0(n4204), .I1(n4205), .S(n4906), .ZN(vectorData1[157])
         );
  MUX4ND0BWP U6273 ( .I0(\vrf/regTable[0][157] ), .I1(\vrf/regTable[1][157] ), 
        .I2(\vrf/regTable[2][157] ), .I3(\vrf/regTable[3][157] ), .S0(n4779), 
        .S1(n4849), .ZN(n4204) );
  MUX4ND0BWP U6274 ( .I0(\vrf/regTable[4][157] ), .I1(\vrf/regTable[5][157] ), 
        .I2(\vrf/regTable[6][157] ), .I3(\vrf/regTable[7][157] ), .S0(n4779), 
        .S1(n4849), .ZN(n4205) );
  MUX2ND0BWP U6275 ( .I0(n4206), .I1(n4207), .S(n4900), .ZN(vectorData1[92])
         );
  MUX4ND0BWP U6276 ( .I0(\vrf/regTable[0][92] ), .I1(\vrf/regTable[1][92] ), 
        .I2(\vrf/regTable[2][92] ), .I3(\vrf/regTable[3][92] ), .S0(n4768), 
        .S1(n4838), .ZN(n4206) );
  MUX4ND0BWP U6277 ( .I0(\vrf/regTable[4][92] ), .I1(\vrf/regTable[5][92] ), 
        .I2(\vrf/regTable[6][92] ), .I3(\vrf/regTable[7][92] ), .S0(n4768), 
        .S1(n4838), .ZN(n4207) );
  MUX2ND0BWP U6278 ( .I0(n4208), .I1(n4209), .S(n4895), .ZN(vectorData1[28])
         );
  MUX4ND0BWP U6279 ( .I0(\vrf/regTable[0][28] ), .I1(\vrf/regTable[1][28] ), 
        .I2(\vrf/regTable[2][28] ), .I3(\vrf/regTable[3][28] ), .S0(n4757), 
        .S1(n4827), .ZN(n4208) );
  MUX4ND0BWP U6280 ( .I0(\vrf/regTable[4][28] ), .I1(\vrf/regTable[5][28] ), 
        .I2(\vrf/regTable[6][28] ), .I3(\vrf/regTable[7][28] ), .S0(n4757), 
        .S1(n4827), .ZN(n4209) );
  MUX2ND0BWP U6281 ( .I0(n4210), .I1(n4211), .S(n4906), .ZN(vectorData1[156])
         );
  MUX4ND0BWP U6282 ( .I0(\vrf/regTable[0][156] ), .I1(\vrf/regTable[1][156] ), 
        .I2(\vrf/regTable[2][156] ), .I3(\vrf/regTable[3][156] ), .S0(n4779), 
        .S1(n4849), .ZN(n4210) );
  MUX4ND0BWP U6283 ( .I0(\vrf/regTable[4][156] ), .I1(\vrf/regTable[5][156] ), 
        .I2(\vrf/regTable[6][156] ), .I3(\vrf/regTable[7][156] ), .S0(n4779), 
        .S1(n4849), .ZN(n4211) );
  MUX2ND0BWP U6284 ( .I0(n4212), .I1(n4213), .S(n4900), .ZN(vectorData1[91])
         );
  MUX4ND0BWP U6285 ( .I0(\vrf/regTable[0][91] ), .I1(\vrf/regTable[1][91] ), 
        .I2(\vrf/regTable[2][91] ), .I3(\vrf/regTable[3][91] ), .S0(n4768), 
        .S1(n4838), .ZN(n4212) );
  MUX4ND0BWP U6286 ( .I0(\vrf/regTable[4][91] ), .I1(\vrf/regTable[5][91] ), 
        .I2(\vrf/regTable[6][91] ), .I3(\vrf/regTable[7][91] ), .S0(n4768), 
        .S1(n4838), .ZN(n4213) );
  MUX2ND0BWP U6287 ( .I0(n4214), .I1(n4215), .S(n4895), .ZN(vectorData1[27])
         );
  MUX4ND0BWP U6288 ( .I0(\vrf/regTable[0][27] ), .I1(\vrf/regTable[1][27] ), 
        .I2(\vrf/regTable[2][27] ), .I3(\vrf/regTable[3][27] ), .S0(n4757), 
        .S1(n4827), .ZN(n4214) );
  MUX4ND0BWP U6289 ( .I0(\vrf/regTable[4][27] ), .I1(\vrf/regTable[5][27] ), 
        .I2(\vrf/regTable[6][27] ), .I3(\vrf/regTable[7][27] ), .S0(n4757), 
        .S1(n4827), .ZN(n4215) );
  MUX2ND0BWP U6290 ( .I0(n4216), .I1(n4217), .S(n4905), .ZN(vectorData1[155])
         );
  MUX4ND0BWP U6291 ( .I0(\vrf/regTable[0][155] ), .I1(\vrf/regTable[1][155] ), 
        .I2(\vrf/regTable[2][155] ), .I3(\vrf/regTable[3][155] ), .S0(n4778), 
        .S1(n4848), .ZN(n4216) );
  MUX4ND0BWP U6292 ( .I0(\vrf/regTable[4][155] ), .I1(\vrf/regTable[5][155] ), 
        .I2(\vrf/regTable[6][155] ), .I3(\vrf/regTable[7][155] ), .S0(n4778), 
        .S1(n4848), .ZN(n4217) );
  MUX2ND0BWP U6293 ( .I0(n4218), .I1(n4219), .S(n4900), .ZN(vectorData1[90])
         );
  MUX4ND0BWP U6294 ( .I0(\vrf/regTable[0][90] ), .I1(\vrf/regTable[1][90] ), 
        .I2(\vrf/regTable[2][90] ), .I3(\vrf/regTable[3][90] ), .S0(n4768), 
        .S1(n4838), .ZN(n4218) );
  MUX4ND0BWP U6295 ( .I0(\vrf/regTable[4][90] ), .I1(\vrf/regTable[5][90] ), 
        .I2(\vrf/regTable[6][90] ), .I3(\vrf/regTable[7][90] ), .S0(n4768), 
        .S1(n4838), .ZN(n4219) );
  MUX2ND0BWP U6296 ( .I0(n4220), .I1(n4221), .S(n4895), .ZN(vectorData1[26])
         );
  MUX4ND0BWP U6297 ( .I0(\vrf/regTable[0][26] ), .I1(\vrf/regTable[1][26] ), 
        .I2(\vrf/regTable[2][26] ), .I3(\vrf/regTable[3][26] ), .S0(n4757), 
        .S1(n4827), .ZN(n4220) );
  MUX4ND0BWP U6298 ( .I0(\vrf/regTable[4][26] ), .I1(\vrf/regTable[5][26] ), 
        .I2(\vrf/regTable[6][26] ), .I3(\vrf/regTable[7][26] ), .S0(n4757), 
        .S1(n4827), .ZN(n4221) );
  MUX2ND0BWP U6299 ( .I0(n4222), .I1(n4223), .S(n4905), .ZN(vectorData1[154])
         );
  MUX4ND0BWP U6300 ( .I0(\vrf/regTable[0][154] ), .I1(\vrf/regTable[1][154] ), 
        .I2(\vrf/regTable[2][154] ), .I3(\vrf/regTable[3][154] ), .S0(n4778), 
        .S1(n4848), .ZN(n4222) );
  MUX4ND0BWP U6301 ( .I0(\vrf/regTable[4][154] ), .I1(\vrf/regTable[5][154] ), 
        .I2(\vrf/regTable[6][154] ), .I3(\vrf/regTable[7][154] ), .S0(n4778), 
        .S1(n4848), .ZN(n4223) );
  MUX2ND0BWP U6302 ( .I0(n4224), .I1(n4225), .S(n4900), .ZN(vectorData1[89])
         );
  MUX4ND0BWP U6303 ( .I0(\vrf/regTable[0][89] ), .I1(\vrf/regTable[1][89] ), 
        .I2(\vrf/regTable[2][89] ), .I3(\vrf/regTable[3][89] ), .S0(n4767), 
        .S1(n4837), .ZN(n4224) );
  MUX4ND0BWP U6304 ( .I0(\vrf/regTable[4][89] ), .I1(\vrf/regTable[5][89] ), 
        .I2(\vrf/regTable[6][89] ), .I3(\vrf/regTable[7][89] ), .S0(n4767), 
        .S1(n4837), .ZN(n4225) );
  MUX2ND0BWP U6305 ( .I0(n4226), .I1(n4227), .S(n4895), .ZN(vectorData1[25])
         );
  MUX4ND0BWP U6306 ( .I0(\vrf/regTable[0][25] ), .I1(\vrf/regTable[1][25] ), 
        .I2(\vrf/regTable[2][25] ), .I3(\vrf/regTable[3][25] ), .S0(n4757), 
        .S1(n4827), .ZN(n4226) );
  MUX4ND0BWP U6307 ( .I0(\vrf/regTable[4][25] ), .I1(\vrf/regTable[5][25] ), 
        .I2(\vrf/regTable[6][25] ), .I3(\vrf/regTable[7][25] ), .S0(n4757), 
        .S1(n4827), .ZN(n4227) );
  MUX2ND0BWP U6308 ( .I0(n4228), .I1(n4229), .S(n4905), .ZN(vectorData1[153])
         );
  MUX4ND0BWP U6309 ( .I0(\vrf/regTable[0][153] ), .I1(\vrf/regTable[1][153] ), 
        .I2(\vrf/regTable[2][153] ), .I3(\vrf/regTable[3][153] ), .S0(n4778), 
        .S1(n4848), .ZN(n4228) );
  MUX4ND0BWP U6310 ( .I0(\vrf/regTable[4][153] ), .I1(\vrf/regTable[5][153] ), 
        .I2(\vrf/regTable[6][153] ), .I3(\vrf/regTable[7][153] ), .S0(n4778), 
        .S1(n4848), .ZN(n4229) );
  MUX2ND0BWP U6311 ( .I0(n4230), .I1(n4231), .S(n4900), .ZN(vectorData1[88])
         );
  MUX4ND0BWP U6312 ( .I0(\vrf/regTable[0][88] ), .I1(\vrf/regTable[1][88] ), 
        .I2(\vrf/regTable[2][88] ), .I3(\vrf/regTable[3][88] ), .S0(n4767), 
        .S1(n4837), .ZN(n4230) );
  MUX4ND0BWP U6313 ( .I0(\vrf/regTable[4][88] ), .I1(\vrf/regTable[5][88] ), 
        .I2(\vrf/regTable[6][88] ), .I3(\vrf/regTable[7][88] ), .S0(n4767), 
        .S1(n4837), .ZN(n4231) );
  MUX2ND0BWP U6314 ( .I0(n4232), .I1(n4233), .S(n4895), .ZN(vectorData1[24])
         );
  MUX4ND0BWP U6315 ( .I0(\vrf/regTable[0][24] ), .I1(\vrf/regTable[1][24] ), 
        .I2(\vrf/regTable[2][24] ), .I3(\vrf/regTable[3][24] ), .S0(n4757), 
        .S1(n4827), .ZN(n4232) );
  MUX4ND0BWP U6316 ( .I0(\vrf/regTable[4][24] ), .I1(\vrf/regTable[5][24] ), 
        .I2(\vrf/regTable[6][24] ), .I3(\vrf/regTable[7][24] ), .S0(n4757), 
        .S1(n4827), .ZN(n4233) );
  MUX2ND0BWP U6317 ( .I0(n4234), .I1(n4235), .S(n4905), .ZN(vectorData1[152])
         );
  MUX4ND0BWP U6318 ( .I0(\vrf/regTable[0][152] ), .I1(\vrf/regTable[1][152] ), 
        .I2(\vrf/regTable[2][152] ), .I3(\vrf/regTable[3][152] ), .S0(n4778), 
        .S1(n4848), .ZN(n4234) );
  MUX4ND0BWP U6319 ( .I0(\vrf/regTable[4][152] ), .I1(\vrf/regTable[5][152] ), 
        .I2(\vrf/regTable[6][152] ), .I3(\vrf/regTable[7][152] ), .S0(n4778), 
        .S1(n4848), .ZN(n4235) );
  MUX2ND0BWP U6320 ( .I0(n4236), .I1(n4237), .S(n4899), .ZN(vectorData1[81])
         );
  MUX4ND0BWP U6321 ( .I0(\vrf/regTable[0][81] ), .I1(\vrf/regTable[1][81] ), 
        .I2(\vrf/regTable[2][81] ), .I3(\vrf/regTable[3][81] ), .S0(n4766), 
        .S1(n4836), .ZN(n4236) );
  MUX4ND0BWP U6322 ( .I0(\vrf/regTable[4][81] ), .I1(\vrf/regTable[5][81] ), 
        .I2(\vrf/regTable[6][81] ), .I3(\vrf/regTable[7][81] ), .S0(n4766), 
        .S1(n4836), .ZN(n4237) );
  MUX2ND0BWP U6323 ( .I0(n4238), .I1(n4239), .S(n4894), .ZN(vectorData1[17])
         );
  MUX4ND0BWP U6324 ( .I0(\vrf/regTable[0][17] ), .I1(\vrf/regTable[1][17] ), 
        .I2(\vrf/regTable[2][17] ), .I3(\vrf/regTable[3][17] ), .S0(n4755), 
        .S1(n4825), .ZN(n4238) );
  MUX4ND0BWP U6325 ( .I0(\vrf/regTable[4][17] ), .I1(\vrf/regTable[5][17] ), 
        .I2(\vrf/regTable[6][17] ), .I3(\vrf/regTable[7][17] ), .S0(n4755), 
        .S1(n4825), .ZN(n4239) );
  MUX2ND0BWP U6326 ( .I0(n4240), .I1(n4241), .S(n4905), .ZN(vectorData1[145])
         );
  MUX4ND0BWP U6327 ( .I0(\vrf/regTable[0][145] ), .I1(\vrf/regTable[1][145] ), 
        .I2(\vrf/regTable[2][145] ), .I3(\vrf/regTable[3][145] ), .S0(n4777), 
        .S1(n4847), .ZN(n4240) );
  MUX4ND0BWP U6328 ( .I0(\vrf/regTable[4][145] ), .I1(\vrf/regTable[5][145] ), 
        .I2(\vrf/regTable[6][145] ), .I3(\vrf/regTable[7][145] ), .S0(n4777), 
        .S1(n4847), .ZN(n4241) );
  MUX2ND0BWP U6329 ( .I0(n4242), .I1(n4243), .S(n4900), .ZN(vectorData1[87])
         );
  MUX4ND0BWP U6330 ( .I0(\vrf/regTable[0][87] ), .I1(\vrf/regTable[1][87] ), 
        .I2(\vrf/regTable[2][87] ), .I3(\vrf/regTable[3][87] ), .S0(n4767), 
        .S1(n4837), .ZN(n4242) );
  MUX4ND0BWP U6331 ( .I0(\vrf/regTable[4][87] ), .I1(\vrf/regTable[5][87] ), 
        .I2(\vrf/regTable[6][87] ), .I3(\vrf/regTable[7][87] ), .S0(n4767), 
        .S1(n4837), .ZN(n4243) );
  MUX2ND0BWP U6332 ( .I0(n4244), .I1(n4245), .S(n4894), .ZN(vectorData1[23])
         );
  MUX4ND0BWP U6333 ( .I0(\vrf/regTable[0][23] ), .I1(\vrf/regTable[1][23] ), 
        .I2(\vrf/regTable[2][23] ), .I3(\vrf/regTable[3][23] ), .S0(n4756), 
        .S1(n4826), .ZN(n4244) );
  MUX4ND0BWP U6334 ( .I0(\vrf/regTable[4][23] ), .I1(\vrf/regTable[5][23] ), 
        .I2(\vrf/regTable[6][23] ), .I3(\vrf/regTable[7][23] ), .S0(n4756), 
        .S1(n4826), .ZN(n4245) );
  MUX2ND0BWP U6335 ( .I0(n4246), .I1(n4247), .S(n4905), .ZN(vectorData1[151])
         );
  MUX4ND0BWP U6336 ( .I0(\vrf/regTable[0][151] ), .I1(\vrf/regTable[1][151] ), 
        .I2(\vrf/regTable[2][151] ), .I3(\vrf/regTable[3][151] ), .S0(n4778), 
        .S1(n4848), .ZN(n4246) );
  MUX4ND0BWP U6337 ( .I0(\vrf/regTable[4][151] ), .I1(\vrf/regTable[5][151] ), 
        .I2(\vrf/regTable[6][151] ), .I3(\vrf/regTable[7][151] ), .S0(n4778), 
        .S1(n4848), .ZN(n4247) );
  MUX2ND0BWP U6338 ( .I0(n4248), .I1(n4249), .S(n4900), .ZN(vectorData1[86])
         );
  MUX4ND0BWP U6339 ( .I0(\vrf/regTable[0][86] ), .I1(\vrf/regTable[1][86] ), 
        .I2(\vrf/regTable[2][86] ), .I3(\vrf/regTable[3][86] ), .S0(n4767), 
        .S1(n4837), .ZN(n4248) );
  MUX4ND0BWP U6340 ( .I0(\vrf/regTable[4][86] ), .I1(\vrf/regTable[5][86] ), 
        .I2(\vrf/regTable[6][86] ), .I3(\vrf/regTable[7][86] ), .S0(n4767), 
        .S1(n4837), .ZN(n4249) );
  MUX2ND0BWP U6341 ( .I0(n4250), .I1(n4251), .S(n4894), .ZN(vectorData1[22])
         );
  MUX4ND0BWP U6342 ( .I0(\vrf/regTable[0][22] ), .I1(\vrf/regTable[1][22] ), 
        .I2(\vrf/regTable[2][22] ), .I3(\vrf/regTable[3][22] ), .S0(n4756), 
        .S1(n4826), .ZN(n4250) );
  MUX4ND0BWP U6343 ( .I0(\vrf/regTable[4][22] ), .I1(\vrf/regTable[5][22] ), 
        .I2(\vrf/regTable[6][22] ), .I3(\vrf/regTable[7][22] ), .S0(n4756), 
        .S1(n4826), .ZN(n4251) );
  MUX2ND0BWP U6344 ( .I0(n4252), .I1(n4253), .S(n4905), .ZN(vectorData1[150])
         );
  MUX4ND0BWP U6345 ( .I0(\vrf/regTable[0][150] ), .I1(\vrf/regTable[1][150] ), 
        .I2(\vrf/regTable[2][150] ), .I3(\vrf/regTable[3][150] ), .S0(n4778), 
        .S1(n4848), .ZN(n4252) );
  MUX4ND0BWP U6346 ( .I0(\vrf/regTable[4][150] ), .I1(\vrf/regTable[5][150] ), 
        .I2(\vrf/regTable[6][150] ), .I3(\vrf/regTable[7][150] ), .S0(n4778), 
        .S1(n4848), .ZN(n4253) );
  MUX2ND0BWP U6347 ( .I0(n4254), .I1(n4255), .S(n4900), .ZN(vectorData1[85])
         );
  MUX4ND0BWP U6348 ( .I0(\vrf/regTable[0][85] ), .I1(\vrf/regTable[1][85] ), 
        .I2(\vrf/regTable[2][85] ), .I3(\vrf/regTable[3][85] ), .S0(n4767), 
        .S1(n4837), .ZN(n4254) );
  MUX4ND0BWP U6349 ( .I0(\vrf/regTable[4][85] ), .I1(\vrf/regTable[5][85] ), 
        .I2(\vrf/regTable[6][85] ), .I3(\vrf/regTable[7][85] ), .S0(n4767), 
        .S1(n4837), .ZN(n4255) );
  MUX2ND0BWP U6350 ( .I0(n4256), .I1(n4257), .S(n4894), .ZN(vectorData1[21])
         );
  MUX4ND0BWP U6351 ( .I0(\vrf/regTable[0][21] ), .I1(\vrf/regTable[1][21] ), 
        .I2(\vrf/regTable[2][21] ), .I3(\vrf/regTable[3][21] ), .S0(n4756), 
        .S1(n4826), .ZN(n4256) );
  MUX4ND0BWP U6352 ( .I0(\vrf/regTable[4][21] ), .I1(\vrf/regTable[5][21] ), 
        .I2(\vrf/regTable[6][21] ), .I3(\vrf/regTable[7][21] ), .S0(n4756), 
        .S1(n4826), .ZN(n4257) );
  MUX2ND0BWP U6353 ( .I0(n4258), .I1(n4259), .S(n4905), .ZN(vectorData1[149])
         );
  MUX4ND0BWP U6354 ( .I0(\vrf/regTable[0][149] ), .I1(\vrf/regTable[1][149] ), 
        .I2(\vrf/regTable[2][149] ), .I3(\vrf/regTable[3][149] ), .S0(n4777), 
        .S1(n4847), .ZN(n4258) );
  MUX4ND0BWP U6355 ( .I0(\vrf/regTable[4][149] ), .I1(\vrf/regTable[5][149] ), 
        .I2(\vrf/regTable[6][149] ), .I3(\vrf/regTable[7][149] ), .S0(n4777), 
        .S1(n4847), .ZN(n4259) );
  MUX2ND0BWP U6356 ( .I0(n4260), .I1(n4261), .S(n4899), .ZN(vectorData1[82])
         );
  MUX4ND0BWP U6357 ( .I0(\vrf/regTable[0][82] ), .I1(\vrf/regTable[1][82] ), 
        .I2(\vrf/regTable[2][82] ), .I3(\vrf/regTable[3][82] ), .S0(n4766), 
        .S1(n4836), .ZN(n4260) );
  MUX4ND0BWP U6358 ( .I0(\vrf/regTable[4][82] ), .I1(\vrf/regTable[5][82] ), 
        .I2(\vrf/regTable[6][82] ), .I3(\vrf/regTable[7][82] ), .S0(n4766), 
        .S1(n4836), .ZN(n4261) );
  MUX2ND0BWP U6359 ( .I0(n4262), .I1(n4263), .S(n4894), .ZN(vectorData1[18])
         );
  MUX4ND0BWP U6360 ( .I0(\vrf/regTable[0][18] ), .I1(\vrf/regTable[1][18] ), 
        .I2(\vrf/regTable[2][18] ), .I3(\vrf/regTable[3][18] ), .S0(n4756), 
        .S1(n4826), .ZN(n4262) );
  MUX4ND0BWP U6361 ( .I0(\vrf/regTable[4][18] ), .I1(\vrf/regTable[5][18] ), 
        .I2(\vrf/regTable[6][18] ), .I3(\vrf/regTable[7][18] ), .S0(n4756), 
        .S1(n4826), .ZN(n4263) );
  MUX2ND0BWP U6362 ( .I0(n4264), .I1(n4265), .S(n4905), .ZN(vectorData1[146])
         );
  MUX4ND0BWP U6363 ( .I0(\vrf/regTable[0][146] ), .I1(\vrf/regTable[1][146] ), 
        .I2(\vrf/regTable[2][146] ), .I3(\vrf/regTable[3][146] ), .S0(n4777), 
        .S1(n4847), .ZN(n4264) );
  MUX4ND0BWP U6364 ( .I0(\vrf/regTable[4][146] ), .I1(\vrf/regTable[5][146] ), 
        .I2(\vrf/regTable[6][146] ), .I3(\vrf/regTable[7][146] ), .S0(n4777), 
        .S1(n4847), .ZN(n4265) );
  MUX2ND0BWP U6365 ( .I0(n4266), .I1(n4267), .S(n4899), .ZN(vectorData1[83])
         );
  MUX4ND0BWP U6366 ( .I0(\vrf/regTable[0][83] ), .I1(\vrf/regTable[1][83] ), 
        .I2(\vrf/regTable[2][83] ), .I3(\vrf/regTable[3][83] ), .S0(n4766), 
        .S1(n4836), .ZN(n4266) );
  MUX4ND0BWP U6367 ( .I0(\vrf/regTable[4][83] ), .I1(\vrf/regTable[5][83] ), 
        .I2(\vrf/regTable[6][83] ), .I3(\vrf/regTable[7][83] ), .S0(n4766), 
        .S1(n4836), .ZN(n4267) );
  MUX2ND0BWP U6368 ( .I0(n4268), .I1(n4269), .S(n4894), .ZN(vectorData1[19])
         );
  MUX4ND0BWP U6369 ( .I0(\vrf/regTable[0][19] ), .I1(\vrf/regTable[1][19] ), 
        .I2(\vrf/regTable[2][19] ), .I3(\vrf/regTable[3][19] ), .S0(n4756), 
        .S1(n4826), .ZN(n4268) );
  MUX4ND0BWP U6370 ( .I0(\vrf/regTable[4][19] ), .I1(\vrf/regTable[5][19] ), 
        .I2(\vrf/regTable[6][19] ), .I3(\vrf/regTable[7][19] ), .S0(n4756), 
        .S1(n4826), .ZN(n4269) );
  MUX2ND0BWP U6371 ( .I0(n4270), .I1(n4271), .S(n4905), .ZN(vectorData1[147])
         );
  MUX4ND0BWP U6372 ( .I0(\vrf/regTable[0][147] ), .I1(\vrf/regTable[1][147] ), 
        .I2(\vrf/regTable[2][147] ), .I3(\vrf/regTable[3][147] ), .S0(n4777), 
        .S1(n4847), .ZN(n4270) );
  MUX4ND0BWP U6373 ( .I0(\vrf/regTable[4][147] ), .I1(\vrf/regTable[5][147] ), 
        .I2(\vrf/regTable[6][147] ), .I3(\vrf/regTable[7][147] ), .S0(n4777), 
        .S1(n4847), .ZN(n4271) );
  MUX2ND0BWP U6374 ( .I0(n4272), .I1(n4273), .S(n4900), .ZN(vectorData1[84])
         );
  MUX4ND0BWP U6375 ( .I0(\vrf/regTable[0][84] ), .I1(\vrf/regTable[1][84] ), 
        .I2(\vrf/regTable[2][84] ), .I3(\vrf/regTable[3][84] ), .S0(n4767), 
        .S1(n4837), .ZN(n4272) );
  MUX4ND0BWP U6376 ( .I0(\vrf/regTable[4][84] ), .I1(\vrf/regTable[5][84] ), 
        .I2(\vrf/regTable[6][84] ), .I3(\vrf/regTable[7][84] ), .S0(n4767), 
        .S1(n4837), .ZN(n4273) );
  MUX2ND0BWP U6377 ( .I0(n4274), .I1(n4275), .S(n4894), .ZN(vectorData1[20])
         );
  MUX4ND0BWP U6378 ( .I0(\vrf/regTable[0][20] ), .I1(\vrf/regTable[1][20] ), 
        .I2(\vrf/regTable[2][20] ), .I3(\vrf/regTable[3][20] ), .S0(n4756), 
        .S1(n4826), .ZN(n4274) );
  MUX4ND0BWP U6379 ( .I0(\vrf/regTable[4][20] ), .I1(\vrf/regTable[5][20] ), 
        .I2(\vrf/regTable[6][20] ), .I3(\vrf/regTable[7][20] ), .S0(n4756), 
        .S1(n4826), .ZN(n4275) );
  MUX2ND0BWP U6380 ( .I0(n4276), .I1(n4277), .S(n4905), .ZN(vectorData1[148])
         );
  MUX4ND0BWP U6381 ( .I0(\vrf/regTable[0][148] ), .I1(\vrf/regTable[1][148] ), 
        .I2(\vrf/regTable[2][148] ), .I3(\vrf/regTable[3][148] ), .S0(n4777), 
        .S1(n4847), .ZN(n4276) );
  MUX4ND0BWP U6382 ( .I0(\vrf/regTable[4][148] ), .I1(\vrf/regTable[5][148] ), 
        .I2(\vrf/regTable[6][148] ), .I3(\vrf/regTable[7][148] ), .S0(n4777), 
        .S1(n4847), .ZN(n4277) );
  MUX2ND0BWP U6383 ( .I0(n4278), .I1(n4279), .S(n5089), .ZN(scalarData2[3]) );
  MUX4ND0BWP U6384 ( .I0(\srf/regTable[0][3] ), .I1(\srf/regTable[1][3] ), 
        .I2(\srf/regTable[2][3] ), .I3(\srf/regTable[3][3] ), .S0(n4971), .S1(
        n5041), .ZN(n4278) );
  MUX4ND0BWP U6385 ( .I0(\srf/regTable[4][3] ), .I1(\srf/regTable[5][3] ), 
        .I2(\srf/regTable[6][3] ), .I3(\srf/regTable[7][3] ), .S0(n4971), .S1(
        n5041), .ZN(n4279) );
  MUX2ND0BWP U6386 ( .I0(n4280), .I1(n4281), .S(n5089), .ZN(scalarData2[4]) );
  MUX4ND0BWP U6387 ( .I0(\srf/regTable[0][4] ), .I1(\srf/regTable[1][4] ), 
        .I2(\srf/regTable[2][4] ), .I3(\srf/regTable[3][4] ), .S0(n4971), .S1(
        n5041), .ZN(n4280) );
  MUX4ND0BWP U6388 ( .I0(\srf/regTable[4][4] ), .I1(\srf/regTable[5][4] ), 
        .I2(\srf/regTable[6][4] ), .I3(\srf/regTable[7][4] ), .S0(n4971), .S1(
        n5041), .ZN(n4281) );
  MUX2ND0BWP U6389 ( .I0(n4282), .I1(n4283), .S(n5074), .ZN(vectorData2[80])
         );
  MUX4ND0BWP U6390 ( .I0(\vrf/regTable[0][80] ), .I1(\vrf/regTable[1][80] ), 
        .I2(\vrf/regTable[2][80] ), .I3(\vrf/regTable[3][80] ), .S0(n4941), 
        .S1(n5011), .ZN(n4282) );
  MUX4ND0BWP U6391 ( .I0(\vrf/regTable[4][80] ), .I1(\vrf/regTable[5][80] ), 
        .I2(\vrf/regTable[6][80] ), .I3(\vrf/regTable[7][80] ), .S0(n4941), 
        .S1(n5011), .ZN(n4283) );
  MUX2ND0BWP U6392 ( .I0(n4284), .I1(n4285), .S(n5074), .ZN(vectorData2[81])
         );
  MUX4ND0BWP U6393 ( .I0(\vrf/regTable[0][81] ), .I1(\vrf/regTable[1][81] ), 
        .I2(\vrf/regTable[2][81] ), .I3(\vrf/regTable[3][81] ), .S0(n4941), 
        .S1(n5011), .ZN(n4284) );
  MUX4ND0BWP U6394 ( .I0(\vrf/regTable[4][81] ), .I1(\vrf/regTable[5][81] ), 
        .I2(\vrf/regTable[6][81] ), .I3(\vrf/regTable[7][81] ), .S0(n4941), 
        .S1(n5011), .ZN(n4285) );
  MUX2ND0BWP U6395 ( .I0(n4286), .I1(n4287), .S(n5075), .ZN(vectorData2[88])
         );
  MUX4ND0BWP U6396 ( .I0(\vrf/regTable[0][88] ), .I1(\vrf/regTable[1][88] ), 
        .I2(\vrf/regTable[2][88] ), .I3(\vrf/regTable[3][88] ), .S0(n4942), 
        .S1(n5012), .ZN(n4286) );
  MUX4ND0BWP U6397 ( .I0(\vrf/regTable[4][88] ), .I1(\vrf/regTable[5][88] ), 
        .I2(\vrf/regTable[6][88] ), .I3(\vrf/regTable[7][88] ), .S0(n4942), 
        .S1(n5012), .ZN(n4287) );
  MUX2ND0BWP U6398 ( .I0(n4288), .I1(n4289), .S(n5075), .ZN(vectorData2[89])
         );
  MUX4ND0BWP U6399 ( .I0(\vrf/regTable[0][89] ), .I1(\vrf/regTable[1][89] ), 
        .I2(\vrf/regTable[2][89] ), .I3(\vrf/regTable[3][89] ), .S0(n4942), 
        .S1(n5012), .ZN(n4288) );
  MUX4ND0BWP U6400 ( .I0(\vrf/regTable[4][89] ), .I1(\vrf/regTable[5][89] ), 
        .I2(\vrf/regTable[6][89] ), .I3(\vrf/regTable[7][89] ), .S0(n4942), 
        .S1(n5012), .ZN(n4289) );
  MUX2ND0BWP U6401 ( .I0(n4290), .I1(n4291), .S(n5075), .ZN(vectorData2[90])
         );
  MUX4ND0BWP U6402 ( .I0(\vrf/regTable[0][90] ), .I1(\vrf/regTable[1][90] ), 
        .I2(\vrf/regTable[2][90] ), .I3(\vrf/regTable[3][90] ), .S0(n4943), 
        .S1(n5013), .ZN(n4290) );
  MUX4ND0BWP U6403 ( .I0(\vrf/regTable[4][90] ), .I1(\vrf/regTable[5][90] ), 
        .I2(\vrf/regTable[6][90] ), .I3(\vrf/regTable[7][90] ), .S0(n4943), 
        .S1(n5013), .ZN(n4291) );
  MUX2ND0BWP U6404 ( .I0(n4292), .I1(n4293), .S(n5075), .ZN(vectorData2[91])
         );
  MUX4ND0BWP U6405 ( .I0(\vrf/regTable[0][91] ), .I1(\vrf/regTable[1][91] ), 
        .I2(\vrf/regTable[2][91] ), .I3(\vrf/regTable[3][91] ), .S0(n4943), 
        .S1(n5013), .ZN(n4292) );
  MUX4ND0BWP U6406 ( .I0(\vrf/regTable[4][91] ), .I1(\vrf/regTable[5][91] ), 
        .I2(\vrf/regTable[6][91] ), .I3(\vrf/regTable[7][91] ), .S0(n4943), 
        .S1(n5013), .ZN(n4293) );
  MUX2ND0BWP U6407 ( .I0(n4294), .I1(n4295), .S(n5075), .ZN(vectorData2[92])
         );
  MUX4ND0BWP U6408 ( .I0(\vrf/regTable[0][92] ), .I1(\vrf/regTable[1][92] ), 
        .I2(\vrf/regTable[2][92] ), .I3(\vrf/regTable[3][92] ), .S0(n4943), 
        .S1(n5013), .ZN(n4294) );
  MUX4ND0BWP U6409 ( .I0(\vrf/regTable[4][92] ), .I1(\vrf/regTable[5][92] ), 
        .I2(\vrf/regTable[6][92] ), .I3(\vrf/regTable[7][92] ), .S0(n4943), 
        .S1(n5013), .ZN(n4295) );
  MUX2ND0BWP U6410 ( .I0(n4296), .I1(n4297), .S(n5075), .ZN(vectorData2[93])
         );
  MUX4ND0BWP U6411 ( .I0(\vrf/regTable[0][93] ), .I1(\vrf/regTable[1][93] ), 
        .I2(\vrf/regTable[2][93] ), .I3(\vrf/regTable[3][93] ), .S0(n4943), 
        .S1(n5013), .ZN(n4296) );
  MUX4ND0BWP U6412 ( .I0(\vrf/regTable[4][93] ), .I1(\vrf/regTable[5][93] ), 
        .I2(\vrf/regTable[6][93] ), .I3(\vrf/regTable[7][93] ), .S0(n4943), 
        .S1(n5013), .ZN(n4297) );
  MUX2ND0BWP U6413 ( .I0(n4298), .I1(n4299), .S(n5075), .ZN(vectorData2[94])
         );
  MUX4ND0BWP U6414 ( .I0(\vrf/regTable[0][94] ), .I1(\vrf/regTable[1][94] ), 
        .I2(\vrf/regTable[2][94] ), .I3(\vrf/regTable[3][94] ), .S0(n4943), 
        .S1(n5013), .ZN(n4298) );
  MUX4ND0BWP U6415 ( .I0(\vrf/regTable[4][94] ), .I1(\vrf/regTable[5][94] ), 
        .I2(\vrf/regTable[6][94] ), .I3(\vrf/regTable[7][94] ), .S0(n4943), 
        .S1(n5013), .ZN(n4299) );
  MUX2ND0BWP U6416 ( .I0(n4300), .I1(n4301), .S(n5075), .ZN(vectorData2[95])
         );
  MUX4ND0BWP U6417 ( .I0(\vrf/regTable[0][95] ), .I1(\vrf/regTable[1][95] ), 
        .I2(\vrf/regTable[2][95] ), .I3(\vrf/regTable[3][95] ), .S0(n4943), 
        .S1(n5013), .ZN(n4300) );
  MUX4ND0BWP U6418 ( .I0(\vrf/regTable[4][95] ), .I1(\vrf/regTable[5][95] ), 
        .I2(\vrf/regTable[6][95] ), .I3(\vrf/regTable[7][95] ), .S0(n4943), 
        .S1(n5013), .ZN(n4301) );
  MUX2ND0BWP U6419 ( .I0(n4302), .I1(n4303), .S(n5074), .ZN(vectorData2[82])
         );
  MUX4ND0BWP U6420 ( .I0(\vrf/regTable[0][82] ), .I1(\vrf/regTable[1][82] ), 
        .I2(\vrf/regTable[2][82] ), .I3(\vrf/regTable[3][82] ), .S0(n4941), 
        .S1(n5011), .ZN(n4302) );
  MUX4ND0BWP U6421 ( .I0(\vrf/regTable[4][82] ), .I1(\vrf/regTable[5][82] ), 
        .I2(\vrf/regTable[6][82] ), .I3(\vrf/regTable[7][82] ), .S0(n4941), 
        .S1(n5011), .ZN(n4303) );
  MUX2ND0BWP U6422 ( .I0(n4304), .I1(n4305), .S(n5075), .ZN(vectorData2[85])
         );
  MUX4ND0BWP U6423 ( .I0(\vrf/regTable[0][85] ), .I1(\vrf/regTable[1][85] ), 
        .I2(\vrf/regTable[2][85] ), .I3(\vrf/regTable[3][85] ), .S0(n4942), 
        .S1(n5012), .ZN(n4304) );
  MUX4ND0BWP U6424 ( .I0(\vrf/regTable[4][85] ), .I1(\vrf/regTable[5][85] ), 
        .I2(\vrf/regTable[6][85] ), .I3(\vrf/regTable[7][85] ), .S0(n4942), 
        .S1(n5012), .ZN(n4305) );
  MUX2ND0BWP U6425 ( .I0(n4306), .I1(n4307), .S(n5075), .ZN(vectorData2[86])
         );
  MUX4ND0BWP U6426 ( .I0(\vrf/regTable[0][86] ), .I1(\vrf/regTable[1][86] ), 
        .I2(\vrf/regTable[2][86] ), .I3(\vrf/regTable[3][86] ), .S0(n4942), 
        .S1(n5012), .ZN(n4306) );
  MUX4ND0BWP U6427 ( .I0(\vrf/regTable[4][86] ), .I1(\vrf/regTable[5][86] ), 
        .I2(\vrf/regTable[6][86] ), .I3(\vrf/regTable[7][86] ), .S0(n4942), 
        .S1(n5012), .ZN(n4307) );
  MUX2ND0BWP U6428 ( .I0(n4308), .I1(n4309), .S(n5075), .ZN(vectorData2[87])
         );
  MUX4ND0BWP U6429 ( .I0(\vrf/regTable[0][87] ), .I1(\vrf/regTable[1][87] ), 
        .I2(\vrf/regTable[2][87] ), .I3(\vrf/regTable[3][87] ), .S0(n4942), 
        .S1(n5012), .ZN(n4308) );
  MUX4ND0BWP U6430 ( .I0(\vrf/regTable[4][87] ), .I1(\vrf/regTable[5][87] ), 
        .I2(\vrf/regTable[6][87] ), .I3(\vrf/regTable[7][87] ), .S0(n4942), 
        .S1(n5012), .ZN(n4309) );
  MUX2ND0BWP U6431 ( .I0(n4310), .I1(n4311), .S(n5085), .ZN(vectorData2[208])
         );
  MUX4ND0BWP U6432 ( .I0(\vrf/regTable[0][208] ), .I1(\vrf/regTable[1][208] ), 
        .I2(\vrf/regTable[2][208] ), .I3(\vrf/regTable[3][208] ), .S0(n4962), 
        .S1(n5032), .ZN(n4310) );
  MUX4ND0BWP U6433 ( .I0(\vrf/regTable[4][208] ), .I1(\vrf/regTable[5][208] ), 
        .I2(\vrf/regTable[6][208] ), .I3(\vrf/regTable[7][208] ), .S0(n4962), 
        .S1(n5032), .ZN(n4311) );
  MUX2ND0BWP U6434 ( .I0(n4312), .I1(n4313), .S(n5081), .ZN(vectorData2[160])
         );
  MUX4ND0BWP U6435 ( .I0(\vrf/regTable[0][160] ), .I1(\vrf/regTable[1][160] ), 
        .I2(\vrf/regTable[2][160] ), .I3(\vrf/regTable[3][160] ), .S0(n4954), 
        .S1(n5024), .ZN(n4312) );
  MUX4ND0BWP U6436 ( .I0(\vrf/regTable[4][160] ), .I1(\vrf/regTable[5][160] ), 
        .I2(\vrf/regTable[6][160] ), .I3(\vrf/regTable[7][160] ), .S0(n4954), 
        .S1(n5024), .ZN(n4313) );
  MUX2ND0BWP U6437 ( .I0(n4314), .I1(n4315), .S(n5072), .ZN(vectorData2[48])
         );
  MUX4ND0BWP U6438 ( .I0(\vrf/regTable[0][48] ), .I1(\vrf/regTable[1][48] ), 
        .I2(\vrf/regTable[2][48] ), .I3(\vrf/regTable[3][48] ), .S0(n4936), 
        .S1(n5006), .ZN(n4314) );
  MUX4ND0BWP U6439 ( .I0(\vrf/regTable[4][48] ), .I1(\vrf/regTable[5][48] ), 
        .I2(\vrf/regTable[6][48] ), .I3(\vrf/regTable[7][48] ), .S0(n4936), 
        .S1(n5006), .ZN(n4315) );
  MUX2ND0BWP U6440 ( .I0(n4316), .I1(n4317), .S(n5085), .ZN(vectorData2[209])
         );
  MUX4ND0BWP U6441 ( .I0(\vrf/regTable[0][209] ), .I1(\vrf/regTable[1][209] ), 
        .I2(\vrf/regTable[2][209] ), .I3(\vrf/regTable[3][209] ), .S0(n4962), 
        .S1(n5032), .ZN(n4316) );
  MUX4ND0BWP U6442 ( .I0(\vrf/regTable[4][209] ), .I1(\vrf/regTable[5][209] ), 
        .I2(\vrf/regTable[6][209] ), .I3(\vrf/regTable[7][209] ), .S0(n4962), 
        .S1(n5032), .ZN(n4317) );
  MUX2ND0BWP U6443 ( .I0(n4318), .I1(n4319), .S(n5081), .ZN(vectorData2[161])
         );
  MUX4ND0BWP U6444 ( .I0(\vrf/regTable[0][161] ), .I1(\vrf/regTable[1][161] ), 
        .I2(\vrf/regTable[2][161] ), .I3(\vrf/regTable[3][161] ), .S0(n4954), 
        .S1(n5024), .ZN(n4318) );
  MUX4ND0BWP U6445 ( .I0(\vrf/regTable[4][161] ), .I1(\vrf/regTable[5][161] ), 
        .I2(\vrf/regTable[6][161] ), .I3(\vrf/regTable[7][161] ), .S0(n4954), 
        .S1(n5024), .ZN(n4319) );
  MUX2ND0BWP U6446 ( .I0(n4320), .I1(n4321), .S(n5072), .ZN(vectorData2[49])
         );
  MUX4ND0BWP U6447 ( .I0(\vrf/regTable[0][49] ), .I1(\vrf/regTable[1][49] ), 
        .I2(\vrf/regTable[2][49] ), .I3(\vrf/regTable[3][49] ), .S0(n4936), 
        .S1(n5006), .ZN(n4320) );
  MUX4ND0BWP U6448 ( .I0(\vrf/regTable[4][49] ), .I1(\vrf/regTable[5][49] ), 
        .I2(\vrf/regTable[6][49] ), .I3(\vrf/regTable[7][49] ), .S0(n4936), 
        .S1(n5006), .ZN(n4321) );
  MUX2ND0BWP U6449 ( .I0(n4322), .I1(n4323), .S(n5086), .ZN(vectorData2[216])
         );
  MUX4ND0BWP U6450 ( .I0(\vrf/regTable[0][216] ), .I1(\vrf/regTable[1][216] ), 
        .I2(\vrf/regTable[2][216] ), .I3(\vrf/regTable[3][216] ), .S0(n4964), 
        .S1(n5034), .ZN(n4322) );
  MUX4ND0BWP U6451 ( .I0(\vrf/regTable[4][216] ), .I1(\vrf/regTable[5][216] ), 
        .I2(\vrf/regTable[6][216] ), .I3(\vrf/regTable[7][216] ), .S0(n4964), 
        .S1(n5034), .ZN(n4323) );
  MUX2ND0BWP U6452 ( .I0(n4324), .I1(n4325), .S(n5082), .ZN(vectorData2[168])
         );
  MUX4ND0BWP U6453 ( .I0(\vrf/regTable[0][168] ), .I1(\vrf/regTable[1][168] ), 
        .I2(\vrf/regTable[2][168] ), .I3(\vrf/regTable[3][168] ), .S0(n4956), 
        .S1(n5026), .ZN(n4324) );
  MUX4ND0BWP U6454 ( .I0(\vrf/regTable[4][168] ), .I1(\vrf/regTable[5][168] ), 
        .I2(\vrf/regTable[6][168] ), .I3(\vrf/regTable[7][168] ), .S0(n4956), 
        .S1(n5026), .ZN(n4325) );
  MUX2ND0BWP U6455 ( .I0(n4326), .I1(n4327), .S(n5072), .ZN(vectorData2[56])
         );
  MUX4ND0BWP U6456 ( .I0(\vrf/regTable[0][56] ), .I1(\vrf/regTable[1][56] ), 
        .I2(\vrf/regTable[2][56] ), .I3(\vrf/regTable[3][56] ), .S0(n4937), 
        .S1(n5007), .ZN(n4326) );
  MUX4ND0BWP U6457 ( .I0(\vrf/regTable[4][56] ), .I1(\vrf/regTable[5][56] ), 
        .I2(\vrf/regTable[6][56] ), .I3(\vrf/regTable[7][56] ), .S0(n4937), 
        .S1(n5007), .ZN(n4327) );
  MUX2ND0BWP U6458 ( .I0(n4328), .I1(n4329), .S(n5086), .ZN(vectorData2[217])
         );
  MUX4ND0BWP U6459 ( .I0(\vrf/regTable[0][217] ), .I1(\vrf/regTable[1][217] ), 
        .I2(\vrf/regTable[2][217] ), .I3(\vrf/regTable[3][217] ), .S0(n4964), 
        .S1(n5034), .ZN(n4328) );
  MUX4ND0BWP U6460 ( .I0(\vrf/regTable[4][217] ), .I1(\vrf/regTable[5][217] ), 
        .I2(\vrf/regTable[6][217] ), .I3(\vrf/regTable[7][217] ), .S0(n4964), 
        .S1(n5034), .ZN(n4329) );
  MUX2ND0BWP U6461 ( .I0(n4330), .I1(n4331), .S(n5082), .ZN(vectorData2[169])
         );
  MUX4ND0BWP U6462 ( .I0(\vrf/regTable[0][169] ), .I1(\vrf/regTable[1][169] ), 
        .I2(\vrf/regTable[2][169] ), .I3(\vrf/regTable[3][169] ), .S0(n4956), 
        .S1(n5026), .ZN(n4330) );
  MUX4ND0BWP U6463 ( .I0(\vrf/regTable[4][169] ), .I1(\vrf/regTable[5][169] ), 
        .I2(\vrf/regTable[6][169] ), .I3(\vrf/regTable[7][169] ), .S0(n4956), 
        .S1(n5026), .ZN(n4331) );
  MUX2ND0BWP U6464 ( .I0(n4332), .I1(n4333), .S(n5072), .ZN(vectorData2[57])
         );
  MUX4ND0BWP U6465 ( .I0(\vrf/regTable[0][57] ), .I1(\vrf/regTable[1][57] ), 
        .I2(\vrf/regTable[2][57] ), .I3(\vrf/regTable[3][57] ), .S0(n4937), 
        .S1(n5007), .ZN(n4332) );
  MUX4ND0BWP U6466 ( .I0(\vrf/regTable[4][57] ), .I1(\vrf/regTable[5][57] ), 
        .I2(\vrf/regTable[6][57] ), .I3(\vrf/regTable[7][57] ), .S0(n4937), 
        .S1(n5007), .ZN(n4333) );
  MUX2ND0BWP U6467 ( .I0(n4334), .I1(n4335), .S(n5086), .ZN(vectorData2[218])
         );
  MUX4ND0BWP U6468 ( .I0(\vrf/regTable[0][218] ), .I1(\vrf/regTable[1][218] ), 
        .I2(\vrf/regTable[2][218] ), .I3(\vrf/regTable[3][218] ), .S0(n4964), 
        .S1(n5034), .ZN(n4334) );
  MUX4ND0BWP U6469 ( .I0(\vrf/regTable[4][218] ), .I1(\vrf/regTable[5][218] ), 
        .I2(\vrf/regTable[6][218] ), .I3(\vrf/regTable[7][218] ), .S0(n4964), 
        .S1(n5034), .ZN(n4335) );
  MUX2ND0BWP U6470 ( .I0(n4336), .I1(n4337), .S(n5082), .ZN(vectorData2[170])
         );
  MUX4ND0BWP U6471 ( .I0(\vrf/regTable[0][170] ), .I1(\vrf/regTable[1][170] ), 
        .I2(\vrf/regTable[2][170] ), .I3(\vrf/regTable[3][170] ), .S0(n4956), 
        .S1(n5026), .ZN(n4336) );
  MUX4ND0BWP U6472 ( .I0(\vrf/regTable[4][170] ), .I1(\vrf/regTable[5][170] ), 
        .I2(\vrf/regTable[6][170] ), .I3(\vrf/regTable[7][170] ), .S0(n4956), 
        .S1(n5026), .ZN(n4337) );
  MUX2ND0BWP U6473 ( .I0(n4338), .I1(n4339), .S(n5072), .ZN(vectorData2[58])
         );
  MUX4ND0BWP U6474 ( .I0(\vrf/regTable[0][58] ), .I1(\vrf/regTable[1][58] ), 
        .I2(\vrf/regTable[2][58] ), .I3(\vrf/regTable[3][58] ), .S0(n4937), 
        .S1(n5007), .ZN(n4338) );
  MUX4ND0BWP U6475 ( .I0(\vrf/regTable[4][58] ), .I1(\vrf/regTable[5][58] ), 
        .I2(\vrf/regTable[6][58] ), .I3(\vrf/regTable[7][58] ), .S0(n4937), 
        .S1(n5007), .ZN(n4339) );
  MUX2ND0BWP U6476 ( .I0(n4340), .I1(n4341), .S(n5086), .ZN(vectorData2[219])
         );
  MUX4ND0BWP U6477 ( .I0(\vrf/regTable[0][219] ), .I1(\vrf/regTable[1][219] ), 
        .I2(\vrf/regTable[2][219] ), .I3(\vrf/regTable[3][219] ), .S0(n4964), 
        .S1(n5034), .ZN(n4340) );
  MUX4ND0BWP U6478 ( .I0(\vrf/regTable[4][219] ), .I1(\vrf/regTable[5][219] ), 
        .I2(\vrf/regTable[6][219] ), .I3(\vrf/regTable[7][219] ), .S0(n4964), 
        .S1(n5034), .ZN(n4341) );
  MUX2ND0BWP U6479 ( .I0(n4342), .I1(n4343), .S(n5082), .ZN(vectorData2[171])
         );
  MUX4ND0BWP U6480 ( .I0(\vrf/regTable[0][171] ), .I1(\vrf/regTable[1][171] ), 
        .I2(\vrf/regTable[2][171] ), .I3(\vrf/regTable[3][171] ), .S0(n4956), 
        .S1(n5026), .ZN(n4342) );
  MUX4ND0BWP U6481 ( .I0(\vrf/regTable[4][171] ), .I1(\vrf/regTable[5][171] ), 
        .I2(\vrf/regTable[6][171] ), .I3(\vrf/regTable[7][171] ), .S0(n4956), 
        .S1(n5026), .ZN(n4343) );
  MUX2ND0BWP U6482 ( .I0(n4344), .I1(n4345), .S(n5072), .ZN(vectorData2[59])
         );
  MUX4ND0BWP U6483 ( .I0(\vrf/regTable[0][59] ), .I1(\vrf/regTable[1][59] ), 
        .I2(\vrf/regTable[2][59] ), .I3(\vrf/regTable[3][59] ), .S0(n4937), 
        .S1(n5007), .ZN(n4344) );
  MUX4ND0BWP U6484 ( .I0(\vrf/regTable[4][59] ), .I1(\vrf/regTable[5][59] ), 
        .I2(\vrf/regTable[6][59] ), .I3(\vrf/regTable[7][59] ), .S0(n4937), 
        .S1(n5007), .ZN(n4345) );
  MUX2ND0BWP U6485 ( .I0(n4346), .I1(n4347), .S(n5086), .ZN(vectorData2[220])
         );
  MUX4ND0BWP U6486 ( .I0(\vrf/regTable[0][220] ), .I1(\vrf/regTable[1][220] ), 
        .I2(\vrf/regTable[2][220] ), .I3(\vrf/regTable[3][220] ), .S0(n4964), 
        .S1(n5034), .ZN(n4346) );
  MUX4ND0BWP U6487 ( .I0(\vrf/regTable[4][220] ), .I1(\vrf/regTable[5][220] ), 
        .I2(\vrf/regTable[6][220] ), .I3(\vrf/regTable[7][220] ), .S0(n4964), 
        .S1(n5034), .ZN(n4347) );
  MUX2ND0BWP U6488 ( .I0(n4348), .I1(n4349), .S(n5082), .ZN(vectorData2[172])
         );
  MUX4ND0BWP U6489 ( .I0(\vrf/regTable[0][172] ), .I1(\vrf/regTable[1][172] ), 
        .I2(\vrf/regTable[2][172] ), .I3(\vrf/regTable[3][172] ), .S0(n4956), 
        .S1(n5026), .ZN(n4348) );
  MUX4ND0BWP U6490 ( .I0(\vrf/regTable[4][172] ), .I1(\vrf/regTable[5][172] ), 
        .I2(\vrf/regTable[6][172] ), .I3(\vrf/regTable[7][172] ), .S0(n4956), 
        .S1(n5026), .ZN(n4349) );
  MUX2ND0BWP U6491 ( .I0(n4350), .I1(n4351), .S(n5073), .ZN(vectorData2[60])
         );
  MUX4ND0BWP U6492 ( .I0(\vrf/regTable[0][60] ), .I1(\vrf/regTable[1][60] ), 
        .I2(\vrf/regTable[2][60] ), .I3(\vrf/regTable[3][60] ), .S0(n4938), 
        .S1(n5008), .ZN(n4350) );
  MUX4ND0BWP U6493 ( .I0(\vrf/regTable[4][60] ), .I1(\vrf/regTable[5][60] ), 
        .I2(\vrf/regTable[6][60] ), .I3(\vrf/regTable[7][60] ), .S0(n4938), 
        .S1(n5008), .ZN(n4351) );
  MUX2ND0BWP U6494 ( .I0(n4352), .I1(n4353), .S(n5086), .ZN(vectorData2[221])
         );
  MUX4ND0BWP U6495 ( .I0(\vrf/regTable[0][221] ), .I1(\vrf/regTable[1][221] ), 
        .I2(\vrf/regTable[2][221] ), .I3(\vrf/regTable[3][221] ), .S0(n4964), 
        .S1(n5034), .ZN(n4352) );
  MUX4ND0BWP U6496 ( .I0(\vrf/regTable[4][221] ), .I1(\vrf/regTable[5][221] ), 
        .I2(\vrf/regTable[6][221] ), .I3(\vrf/regTable[7][221] ), .S0(n4964), 
        .S1(n5034), .ZN(n4353) );
  MUX2ND0BWP U6497 ( .I0(n4354), .I1(n4355), .S(n5082), .ZN(vectorData2[173])
         );
  MUX4ND0BWP U6498 ( .I0(\vrf/regTable[0][173] ), .I1(\vrf/regTable[1][173] ), 
        .I2(\vrf/regTable[2][173] ), .I3(\vrf/regTable[3][173] ), .S0(n4956), 
        .S1(n5026), .ZN(n4354) );
  MUX4ND0BWP U6499 ( .I0(\vrf/regTable[4][173] ), .I1(\vrf/regTable[5][173] ), 
        .I2(\vrf/regTable[6][173] ), .I3(\vrf/regTable[7][173] ), .S0(n4956), 
        .S1(n5026), .ZN(n4355) );
  MUX2ND0BWP U6500 ( .I0(n4356), .I1(n4357), .S(n5073), .ZN(vectorData2[61])
         );
  MUX4ND0BWP U6501 ( .I0(\vrf/regTable[0][61] ), .I1(\vrf/regTable[1][61] ), 
        .I2(\vrf/regTable[2][61] ), .I3(\vrf/regTable[3][61] ), .S0(n4938), 
        .S1(n5008), .ZN(n4356) );
  MUX4ND0BWP U6502 ( .I0(\vrf/regTable[4][61] ), .I1(\vrf/regTable[5][61] ), 
        .I2(\vrf/regTable[6][61] ), .I3(\vrf/regTable[7][61] ), .S0(n4938), 
        .S1(n5008), .ZN(n4357) );
  MUX2ND0BWP U6503 ( .I0(n4358), .I1(n4359), .S(n5086), .ZN(vectorData2[222])
         );
  MUX4ND0BWP U6504 ( .I0(\vrf/regTable[0][222] ), .I1(\vrf/regTable[1][222] ), 
        .I2(\vrf/regTable[2][222] ), .I3(\vrf/regTable[3][222] ), .S0(n4965), 
        .S1(n5035), .ZN(n4358) );
  MUX4ND0BWP U6505 ( .I0(\vrf/regTable[4][222] ), .I1(\vrf/regTable[5][222] ), 
        .I2(\vrf/regTable[6][222] ), .I3(\vrf/regTable[7][222] ), .S0(n4965), 
        .S1(n5035), .ZN(n4359) );
  MUX2ND0BWP U6506 ( .I0(n4360), .I1(n4361), .S(n5082), .ZN(vectorData2[174])
         );
  MUX4ND0BWP U6507 ( .I0(\vrf/regTable[0][174] ), .I1(\vrf/regTable[1][174] ), 
        .I2(\vrf/regTable[2][174] ), .I3(\vrf/regTable[3][174] ), .S0(n4957), 
        .S1(n5027), .ZN(n4360) );
  MUX4ND0BWP U6508 ( .I0(\vrf/regTable[4][174] ), .I1(\vrf/regTable[5][174] ), 
        .I2(\vrf/regTable[6][174] ), .I3(\vrf/regTable[7][174] ), .S0(n4957), 
        .S1(n5027), .ZN(n4361) );
  MUX2ND0BWP U6509 ( .I0(n4362), .I1(n4363), .S(n5073), .ZN(vectorData2[62])
         );
  MUX4ND0BWP U6510 ( .I0(\vrf/regTable[0][62] ), .I1(\vrf/regTable[1][62] ), 
        .I2(\vrf/regTable[2][62] ), .I3(\vrf/regTable[3][62] ), .S0(n4938), 
        .S1(n5008), .ZN(n4362) );
  MUX4ND0BWP U6511 ( .I0(\vrf/regTable[4][62] ), .I1(\vrf/regTable[5][62] ), 
        .I2(\vrf/regTable[6][62] ), .I3(\vrf/regTable[7][62] ), .S0(n4938), 
        .S1(n5008), .ZN(n4363) );
  MUX2ND0BWP U6512 ( .I0(n4364), .I1(n4365), .S(n5086), .ZN(vectorData2[223])
         );
  MUX4ND0BWP U6513 ( .I0(\vrf/regTable[0][223] ), .I1(\vrf/regTable[1][223] ), 
        .I2(\vrf/regTable[2][223] ), .I3(\vrf/regTable[3][223] ), .S0(n4965), 
        .S1(n5035), .ZN(n4364) );
  MUX4ND0BWP U6514 ( .I0(\vrf/regTable[4][223] ), .I1(\vrf/regTable[5][223] ), 
        .I2(\vrf/regTable[6][223] ), .I3(\vrf/regTable[7][223] ), .S0(n4965), 
        .S1(n5035), .ZN(n4365) );
  MUX2ND0BWP U6515 ( .I0(n4366), .I1(n4367), .S(n5082), .ZN(vectorData2[175])
         );
  MUX4ND0BWP U6516 ( .I0(\vrf/regTable[0][175] ), .I1(\vrf/regTable[1][175] ), 
        .I2(\vrf/regTable[2][175] ), .I3(\vrf/regTable[3][175] ), .S0(n4957), 
        .S1(n5027), .ZN(n4366) );
  MUX4ND0BWP U6517 ( .I0(\vrf/regTable[4][175] ), .I1(\vrf/regTable[5][175] ), 
        .I2(\vrf/regTable[6][175] ), .I3(\vrf/regTable[7][175] ), .S0(n4957), 
        .S1(n5027), .ZN(n4367) );
  MUX2ND0BWP U6518 ( .I0(n4368), .I1(n4369), .S(n5073), .ZN(vectorData2[63])
         );
  MUX4ND0BWP U6519 ( .I0(\vrf/regTable[0][63] ), .I1(\vrf/regTable[1][63] ), 
        .I2(\vrf/regTable[2][63] ), .I3(\vrf/regTable[3][63] ), .S0(n4938), 
        .S1(n5008), .ZN(n4368) );
  MUX4ND0BWP U6520 ( .I0(\vrf/regTable[4][63] ), .I1(\vrf/regTable[5][63] ), 
        .I2(\vrf/regTable[6][63] ), .I3(\vrf/regTable[7][63] ), .S0(n4938), 
        .S1(n5008), .ZN(n4369) );
  MUX2ND0BWP U6521 ( .I0(n4370), .I1(n4371), .S(n5085), .ZN(vectorData2[210])
         );
  MUX4ND0BWP U6522 ( .I0(\vrf/regTable[0][210] ), .I1(\vrf/regTable[1][210] ), 
        .I2(\vrf/regTable[2][210] ), .I3(\vrf/regTable[3][210] ), .S0(n4963), 
        .S1(n5033), .ZN(n4370) );
  MUX4ND0BWP U6523 ( .I0(\vrf/regTable[4][210] ), .I1(\vrf/regTable[5][210] ), 
        .I2(\vrf/regTable[6][210] ), .I3(\vrf/regTable[7][210] ), .S0(n4963), 
        .S1(n5033), .ZN(n4371) );
  MUX2ND0BWP U6524 ( .I0(n4372), .I1(n4373), .S(n5081), .ZN(vectorData2[162])
         );
  MUX4ND0BWP U6525 ( .I0(\vrf/regTable[0][162] ), .I1(\vrf/regTable[1][162] ), 
        .I2(\vrf/regTable[2][162] ), .I3(\vrf/regTable[3][162] ), .S0(n4955), 
        .S1(n5025), .ZN(n4372) );
  MUX4ND0BWP U6526 ( .I0(\vrf/regTable[4][162] ), .I1(\vrf/regTable[5][162] ), 
        .I2(\vrf/regTable[6][162] ), .I3(\vrf/regTable[7][162] ), .S0(n4955), 
        .S1(n5025), .ZN(n4373) );
  MUX2ND0BWP U6527 ( .I0(n4374), .I1(n4375), .S(n5072), .ZN(vectorData2[50])
         );
  MUX4ND0BWP U6528 ( .I0(\vrf/regTable[0][50] ), .I1(\vrf/regTable[1][50] ), 
        .I2(\vrf/regTable[2][50] ), .I3(\vrf/regTable[3][50] ), .S0(n4936), 
        .S1(n5006), .ZN(n4374) );
  MUX4ND0BWP U6529 ( .I0(\vrf/regTable[4][50] ), .I1(\vrf/regTable[5][50] ), 
        .I2(\vrf/regTable[6][50] ), .I3(\vrf/regTable[7][50] ), .S0(n4936), 
        .S1(n5006), .ZN(n4375) );
  MUX2ND0BWP U6530 ( .I0(n4376), .I1(n4377), .S(n5085), .ZN(vectorData2[213])
         );
  MUX4ND0BWP U6531 ( .I0(\vrf/regTable[0][213] ), .I1(\vrf/regTable[1][213] ), 
        .I2(\vrf/regTable[2][213] ), .I3(\vrf/regTable[3][213] ), .S0(n4963), 
        .S1(n5033), .ZN(n4376) );
  MUX4ND0BWP U6532 ( .I0(\vrf/regTable[4][213] ), .I1(\vrf/regTable[5][213] ), 
        .I2(\vrf/regTable[6][213] ), .I3(\vrf/regTable[7][213] ), .S0(n4963), 
        .S1(n5033), .ZN(n4377) );
  MUX2ND0BWP U6533 ( .I0(n4378), .I1(n4379), .S(n5081), .ZN(vectorData2[165])
         );
  MUX4ND0BWP U6534 ( .I0(\vrf/regTable[0][165] ), .I1(\vrf/regTable[1][165] ), 
        .I2(\vrf/regTable[2][165] ), .I3(\vrf/regTable[3][165] ), .S0(n4955), 
        .S1(n5025), .ZN(n4378) );
  MUX4ND0BWP U6535 ( .I0(\vrf/regTable[4][165] ), .I1(\vrf/regTable[5][165] ), 
        .I2(\vrf/regTable[6][165] ), .I3(\vrf/regTable[7][165] ), .S0(n4955), 
        .S1(n5025), .ZN(n4379) );
  MUX2ND0BWP U6536 ( .I0(n4380), .I1(n4381), .S(n5072), .ZN(vectorData2[53])
         );
  MUX4ND0BWP U6537 ( .I0(\vrf/regTable[0][53] ), .I1(\vrf/regTable[1][53] ), 
        .I2(\vrf/regTable[2][53] ), .I3(\vrf/regTable[3][53] ), .S0(n4936), 
        .S1(n5006), .ZN(n4380) );
  MUX4ND0BWP U6538 ( .I0(\vrf/regTable[4][53] ), .I1(\vrf/regTable[5][53] ), 
        .I2(\vrf/regTable[6][53] ), .I3(\vrf/regTable[7][53] ), .S0(n4936), 
        .S1(n5006), .ZN(n4381) );
  MUX2ND0BWP U6539 ( .I0(n4382), .I1(n4383), .S(n5085), .ZN(vectorData2[214])
         );
  MUX4ND0BWP U6540 ( .I0(\vrf/regTable[0][214] ), .I1(\vrf/regTable[1][214] ), 
        .I2(\vrf/regTable[2][214] ), .I3(\vrf/regTable[3][214] ), .S0(n4963), 
        .S1(n5033), .ZN(n4382) );
  MUX4ND0BWP U6541 ( .I0(\vrf/regTable[4][214] ), .I1(\vrf/regTable[5][214] ), 
        .I2(\vrf/regTable[6][214] ), .I3(\vrf/regTable[7][214] ), .S0(n4963), 
        .S1(n5033), .ZN(n4383) );
  MUX2ND0BWP U6542 ( .I0(n4384), .I1(n4385), .S(n5081), .ZN(vectorData2[166])
         );
  MUX4ND0BWP U6543 ( .I0(\vrf/regTable[0][166] ), .I1(\vrf/regTable[1][166] ), 
        .I2(\vrf/regTable[2][166] ), .I3(\vrf/regTable[3][166] ), .S0(n4955), 
        .S1(n5025), .ZN(n4384) );
  MUX4ND0BWP U6544 ( .I0(\vrf/regTable[4][166] ), .I1(\vrf/regTable[5][166] ), 
        .I2(\vrf/regTable[6][166] ), .I3(\vrf/regTable[7][166] ), .S0(n4955), 
        .S1(n5025), .ZN(n4385) );
  MUX2ND0BWP U6545 ( .I0(n4386), .I1(n4387), .S(n5072), .ZN(vectorData2[54])
         );
  MUX4ND0BWP U6546 ( .I0(\vrf/regTable[0][54] ), .I1(\vrf/regTable[1][54] ), 
        .I2(\vrf/regTable[2][54] ), .I3(\vrf/regTable[3][54] ), .S0(n4937), 
        .S1(n5007), .ZN(n4386) );
  MUX4ND0BWP U6547 ( .I0(\vrf/regTable[4][54] ), .I1(\vrf/regTable[5][54] ), 
        .I2(\vrf/regTable[6][54] ), .I3(\vrf/regTable[7][54] ), .S0(n4937), 
        .S1(n5007), .ZN(n4387) );
  MUX2ND0BWP U6548 ( .I0(n4388), .I1(n4389), .S(n5085), .ZN(vectorData2[215])
         );
  MUX4ND0BWP U6549 ( .I0(\vrf/regTable[0][215] ), .I1(\vrf/regTable[1][215] ), 
        .I2(\vrf/regTable[2][215] ), .I3(\vrf/regTable[3][215] ), .S0(n4963), 
        .S1(n5033), .ZN(n4388) );
  MUX4ND0BWP U6550 ( .I0(\vrf/regTable[4][215] ), .I1(\vrf/regTable[5][215] ), 
        .I2(\vrf/regTable[6][215] ), .I3(\vrf/regTable[7][215] ), .S0(n4963), 
        .S1(n5033), .ZN(n4389) );
  MUX2ND0BWP U6551 ( .I0(n4390), .I1(n4391), .S(n5081), .ZN(vectorData2[167])
         );
  MUX4ND0BWP U6552 ( .I0(\vrf/regTable[0][167] ), .I1(\vrf/regTable[1][167] ), 
        .I2(\vrf/regTable[2][167] ), .I3(\vrf/regTable[3][167] ), .S0(n4955), 
        .S1(n5025), .ZN(n4390) );
  MUX4ND0BWP U6553 ( .I0(\vrf/regTable[4][167] ), .I1(\vrf/regTable[5][167] ), 
        .I2(\vrf/regTable[6][167] ), .I3(\vrf/regTable[7][167] ), .S0(n4955), 
        .S1(n5025), .ZN(n4391) );
  MUX2ND0BWP U6554 ( .I0(n4392), .I1(n4393), .S(n5072), .ZN(vectorData2[55])
         );
  MUX4ND0BWP U6555 ( .I0(\vrf/regTable[0][55] ), .I1(\vrf/regTable[1][55] ), 
        .I2(\vrf/regTable[2][55] ), .I3(\vrf/regTable[3][55] ), .S0(n4937), 
        .S1(n5007), .ZN(n4392) );
  MUX4ND0BWP U6556 ( .I0(\vrf/regTable[4][55] ), .I1(\vrf/regTable[5][55] ), 
        .I2(\vrf/regTable[6][55] ), .I3(\vrf/regTable[7][55] ), .S0(n4937), 
        .S1(n5007), .ZN(n4393) );
  MUX2ND0BWP U6557 ( .I0(n4394), .I1(n4395), .S(n5068), .ZN(vectorData2[3]) );
  MUX4ND0BWP U6558 ( .I0(\vrf/regTable[0][3] ), .I1(\vrf/regTable[1][3] ), 
        .I2(\vrf/regTable[2][3] ), .I3(\vrf/regTable[3][3] ), .S0(n4928), .S1(
        n4998), .ZN(n4394) );
  MUX4ND0BWP U6559 ( .I0(\vrf/regTable[4][3] ), .I1(\vrf/regTable[5][3] ), 
        .I2(\vrf/regTable[6][3] ), .I3(\vrf/regTable[7][3] ), .S0(n4928), .S1(
        n4998), .ZN(n4395) );
  MUX2ND0BWP U6560 ( .I0(n4396), .I1(n4397), .S(n5068), .ZN(vectorData2[4]) );
  MUX4ND0BWP U6561 ( .I0(\vrf/regTable[0][4] ), .I1(\vrf/regTable[1][4] ), 
        .I2(\vrf/regTable[2][4] ), .I3(\vrf/regTable[3][4] ), .S0(n4928), .S1(
        n4998), .ZN(n4396) );
  MUX4ND0BWP U6562 ( .I0(\vrf/regTable[4][4] ), .I1(\vrf/regTable[5][4] ), 
        .I2(\vrf/regTable[6][4] ), .I3(\vrf/regTable[7][4] ), .S0(n4928), .S1(
        n4998), .ZN(n4397) );
  MUX2ND0BWP U6563 ( .I0(n4398), .I1(n4399), .S(n5090), .ZN(scalarData2[11])
         );
  MUX4ND0BWP U6564 ( .I0(\srf/regTable[0][11] ), .I1(\srf/regTable[1][11] ), 
        .I2(\srf/regTable[2][11] ), .I3(\srf/regTable[3][11] ), .S0(n4972), 
        .S1(n5042), .ZN(n4398) );
  MUX4ND0BWP U6565 ( .I0(\srf/regTable[4][11] ), .I1(\srf/regTable[5][11] ), 
        .I2(\srf/regTable[6][11] ), .I3(\srf/regTable[7][11] ), .S0(n4972), 
        .S1(n5042), .ZN(n4399) );
  MUX2ND0BWP U6566 ( .I0(n4400), .I1(n4401), .S(n5090), .ZN(scalarData2[12])
         );
  MUX4ND0BWP U6567 ( .I0(\srf/regTable[0][12] ), .I1(\srf/regTable[1][12] ), 
        .I2(\srf/regTable[2][12] ), .I3(\srf/regTable[3][12] ), .S0(n4972), 
        .S1(n5042), .ZN(n4400) );
  MUX4ND0BWP U6568 ( .I0(\srf/regTable[4][12] ), .I1(\srf/regTable[5][12] ), 
        .I2(\srf/regTable[6][12] ), .I3(\srf/regTable[7][12] ), .S0(n4972), 
        .S1(n5042), .ZN(n4401) );
  MUX2ND0BWP U6569 ( .I0(n4402), .I1(n4403), .S(n5090), .ZN(scalarData2[13])
         );
  MUX4ND0BWP U6570 ( .I0(\srf/regTable[0][13] ), .I1(\srf/regTable[1][13] ), 
        .I2(\srf/regTable[2][13] ), .I3(\srf/regTable[3][13] ), .S0(n4972), 
        .S1(n5042), .ZN(n4402) );
  MUX4ND0BWP U6571 ( .I0(\srf/regTable[4][13] ), .I1(\srf/regTable[5][13] ), 
        .I2(\srf/regTable[6][13] ), .I3(\srf/regTable[7][13] ), .S0(n4972), 
        .S1(n5042), .ZN(n4403) );
  MUX2ND0BWP U6572 ( .I0(n4404), .I1(n4405), .S(n5090), .ZN(scalarData2[14])
         );
  MUX4ND0BWP U6573 ( .I0(\srf/regTable[0][14] ), .I1(\srf/regTable[1][14] ), 
        .I2(\srf/regTable[2][14] ), .I3(\srf/regTable[3][14] ), .S0(n4973), 
        .S1(n5043), .ZN(n4404) );
  MUX4ND0BWP U6574 ( .I0(\srf/regTable[4][14] ), .I1(\srf/regTable[5][14] ), 
        .I2(\srf/regTable[6][14] ), .I3(\srf/regTable[7][14] ), .S0(n4973), 
        .S1(n5043), .ZN(n4405) );
  MUX2ND0BWP U6575 ( .I0(n4406), .I1(n4407), .S(n5090), .ZN(scalarData2[15])
         );
  MUX4ND0BWP U6576 ( .I0(\srf/regTable[0][15] ), .I1(\srf/regTable[1][15] ), 
        .I2(\srf/regTable[2][15] ), .I3(\srf/regTable[3][15] ), .S0(n4973), 
        .S1(n5043), .ZN(n4406) );
  MUX4ND0BWP U6577 ( .I0(\srf/regTable[4][15] ), .I1(\srf/regTable[5][15] ), 
        .I2(\srf/regTable[6][15] ), .I3(\srf/regTable[7][15] ), .S0(n4973), 
        .S1(n5043), .ZN(n4407) );
  MUX2ND0BWP U6578 ( .I0(n4408), .I1(n4409), .S(n5086), .ZN(vectorData2[227])
         );
  MUX4ND0BWP U6579 ( .I0(\vrf/regTable[0][227] ), .I1(\vrf/regTable[1][227] ), 
        .I2(\vrf/regTable[2][227] ), .I3(\vrf/regTable[3][227] ), .S0(n4965), 
        .S1(n5035), .ZN(n4408) );
  MUX4ND0BWP U6580 ( .I0(\vrf/regTable[4][227] ), .I1(\vrf/regTable[5][227] ), 
        .I2(\vrf/regTable[6][227] ), .I3(\vrf/regTable[7][227] ), .S0(n4965), 
        .S1(n5035), .ZN(n4409) );
  MUX2ND0BWP U6581 ( .I0(n4410), .I1(n4411), .S(n5087), .ZN(vectorData2[228])
         );
  MUX4ND0BWP U6582 ( .I0(\vrf/regTable[0][228] ), .I1(\vrf/regTable[1][228] ), 
        .I2(\vrf/regTable[2][228] ), .I3(\vrf/regTable[3][228] ), .S0(n4966), 
        .S1(n5036), .ZN(n4410) );
  MUX4ND0BWP U6583 ( .I0(\vrf/regTable[4][228] ), .I1(\vrf/regTable[5][228] ), 
        .I2(\vrf/regTable[6][228] ), .I3(\vrf/regTable[7][228] ), .S0(n4966), 
        .S1(n5036), .ZN(n4411) );
  MUX2ND0BWP U6584 ( .I0(n4412), .I1(n4413), .S(n5073), .ZN(vectorData2[64])
         );
  MUX4ND0BWP U6585 ( .I0(\vrf/regTable[0][64] ), .I1(\vrf/regTable[1][64] ), 
        .I2(\vrf/regTable[2][64] ), .I3(\vrf/regTable[3][64] ), .S0(n4938), 
        .S1(n5008), .ZN(n4412) );
  MUX4ND0BWP U6586 ( .I0(\vrf/regTable[4][64] ), .I1(\vrf/regTable[5][64] ), 
        .I2(\vrf/regTable[6][64] ), .I3(\vrf/regTable[7][64] ), .S0(n4938), 
        .S1(n5008), .ZN(n4413) );
  MUX2ND0BWP U6587 ( .I0(n4414), .I1(n4415), .S(n5073), .ZN(vectorData2[65])
         );
  MUX4ND0BWP U6588 ( .I0(\vrf/regTable[0][65] ), .I1(\vrf/regTable[1][65] ), 
        .I2(\vrf/regTable[2][65] ), .I3(\vrf/regTable[3][65] ), .S0(n4938), 
        .S1(n5008), .ZN(n4414) );
  MUX4ND0BWP U6589 ( .I0(\vrf/regTable[4][65] ), .I1(\vrf/regTable[5][65] ), 
        .I2(\vrf/regTable[6][65] ), .I3(\vrf/regTable[7][65] ), .S0(n4938), 
        .S1(n5008), .ZN(n4415) );
  MUX2ND0BWP U6590 ( .I0(n4416), .I1(n4417), .S(n5074), .ZN(vectorData2[72])
         );
  MUX4ND0BWP U6591 ( .I0(\vrf/regTable[0][72] ), .I1(\vrf/regTable[1][72] ), 
        .I2(\vrf/regTable[2][72] ), .I3(\vrf/regTable[3][72] ), .S0(n4940), 
        .S1(n5010), .ZN(n4416) );
  MUX4ND0BWP U6592 ( .I0(\vrf/regTable[4][72] ), .I1(\vrf/regTable[5][72] ), 
        .I2(\vrf/regTable[6][72] ), .I3(\vrf/regTable[7][72] ), .S0(n4940), 
        .S1(n5010), .ZN(n4417) );
  MUX2ND0BWP U6593 ( .I0(n4418), .I1(n4419), .S(n5074), .ZN(vectorData2[73])
         );
  MUX4ND0BWP U6594 ( .I0(\vrf/regTable[0][73] ), .I1(\vrf/regTable[1][73] ), 
        .I2(\vrf/regTable[2][73] ), .I3(\vrf/regTable[3][73] ), .S0(n4940), 
        .S1(n5010), .ZN(n4418) );
  MUX4ND0BWP U6595 ( .I0(\vrf/regTable[4][73] ), .I1(\vrf/regTable[5][73] ), 
        .I2(\vrf/regTable[6][73] ), .I3(\vrf/regTable[7][73] ), .S0(n4940), 
        .S1(n5010), .ZN(n4419) );
  MUX2ND0BWP U6596 ( .I0(n4420), .I1(n4421), .S(n5074), .ZN(vectorData2[74])
         );
  MUX4ND0BWP U6597 ( .I0(\vrf/regTable[0][74] ), .I1(\vrf/regTable[1][74] ), 
        .I2(\vrf/regTable[2][74] ), .I3(\vrf/regTable[3][74] ), .S0(n4940), 
        .S1(n5010), .ZN(n4420) );
  MUX4ND0BWP U6598 ( .I0(\vrf/regTable[4][74] ), .I1(\vrf/regTable[5][74] ), 
        .I2(\vrf/regTable[6][74] ), .I3(\vrf/regTable[7][74] ), .S0(n4940), 
        .S1(n5010), .ZN(n4421) );
  MUX2ND0BWP U6599 ( .I0(n4422), .I1(n4423), .S(n5074), .ZN(vectorData2[75])
         );
  MUX4ND0BWP U6600 ( .I0(\vrf/regTable[0][75] ), .I1(\vrf/regTable[1][75] ), 
        .I2(\vrf/regTable[2][75] ), .I3(\vrf/regTable[3][75] ), .S0(n4940), 
        .S1(n5010), .ZN(n4422) );
  MUX4ND0BWP U6601 ( .I0(\vrf/regTable[4][75] ), .I1(\vrf/regTable[5][75] ), 
        .I2(\vrf/regTable[6][75] ), .I3(\vrf/regTable[7][75] ), .S0(n4940), 
        .S1(n5010), .ZN(n4423) );
  MUX2ND0BWP U6602 ( .I0(n4424), .I1(n4425), .S(n5074), .ZN(vectorData2[76])
         );
  MUX4ND0BWP U6603 ( .I0(\vrf/regTable[0][76] ), .I1(\vrf/regTable[1][76] ), 
        .I2(\vrf/regTable[2][76] ), .I3(\vrf/regTable[3][76] ), .S0(n4940), 
        .S1(n5010), .ZN(n4424) );
  MUX4ND0BWP U6604 ( .I0(\vrf/regTable[4][76] ), .I1(\vrf/regTable[5][76] ), 
        .I2(\vrf/regTable[6][76] ), .I3(\vrf/regTable[7][76] ), .S0(n4940), 
        .S1(n5010), .ZN(n4425) );
  MUX2ND0BWP U6605 ( .I0(n4426), .I1(n4427), .S(n5074), .ZN(vectorData2[77])
         );
  MUX4ND0BWP U6606 ( .I0(\vrf/regTable[0][77] ), .I1(\vrf/regTable[1][77] ), 
        .I2(\vrf/regTable[2][77] ), .I3(\vrf/regTable[3][77] ), .S0(n4940), 
        .S1(n5010), .ZN(n4426) );
  MUX4ND0BWP U6607 ( .I0(\vrf/regTable[4][77] ), .I1(\vrf/regTable[5][77] ), 
        .I2(\vrf/regTable[6][77] ), .I3(\vrf/regTable[7][77] ), .S0(n4940), 
        .S1(n5010), .ZN(n4427) );
  MUX2ND0BWP U6608 ( .I0(n4428), .I1(n4429), .S(n5074), .ZN(vectorData2[78])
         );
  MUX4ND0BWP U6609 ( .I0(\vrf/regTable[0][78] ), .I1(\vrf/regTable[1][78] ), 
        .I2(\vrf/regTable[2][78] ), .I3(\vrf/regTable[3][78] ), .S0(n4941), 
        .S1(n5011), .ZN(n4428) );
  MUX4ND0BWP U6610 ( .I0(\vrf/regTable[4][78] ), .I1(\vrf/regTable[5][78] ), 
        .I2(\vrf/regTable[6][78] ), .I3(\vrf/regTable[7][78] ), .S0(n4941), 
        .S1(n5011), .ZN(n4429) );
  MUX2ND0BWP U6611 ( .I0(n4430), .I1(n4431), .S(n5074), .ZN(vectorData2[79])
         );
  MUX4ND0BWP U6612 ( .I0(\vrf/regTable[0][79] ), .I1(\vrf/regTable[1][79] ), 
        .I2(\vrf/regTable[2][79] ), .I3(\vrf/regTable[3][79] ), .S0(n4941), 
        .S1(n5011), .ZN(n4430) );
  MUX4ND0BWP U6613 ( .I0(\vrf/regTable[4][79] ), .I1(\vrf/regTable[5][79] ), 
        .I2(\vrf/regTable[6][79] ), .I3(\vrf/regTable[7][79] ), .S0(n4941), 
        .S1(n5011), .ZN(n4431) );
  MUX2ND0BWP U6614 ( .I0(n4432), .I1(n4433), .S(n5073), .ZN(vectorData2[66])
         );
  MUX4ND0BWP U6615 ( .I0(\vrf/regTable[0][66] ), .I1(\vrf/regTable[1][66] ), 
        .I2(\vrf/regTable[2][66] ), .I3(\vrf/regTable[3][66] ), .S0(n4939), 
        .S1(n5009), .ZN(n4432) );
  MUX4ND0BWP U6616 ( .I0(\vrf/regTable[4][66] ), .I1(\vrf/regTable[5][66] ), 
        .I2(\vrf/regTable[6][66] ), .I3(\vrf/regTable[7][66] ), .S0(n4939), 
        .S1(n5009), .ZN(n4433) );
  MUX2ND0BWP U6617 ( .I0(n4434), .I1(n4435), .S(n5073), .ZN(vectorData2[69])
         );
  MUX4ND0BWP U6618 ( .I0(\vrf/regTable[0][69] ), .I1(\vrf/regTable[1][69] ), 
        .I2(\vrf/regTable[2][69] ), .I3(\vrf/regTable[3][69] ), .S0(n4939), 
        .S1(n5009), .ZN(n4434) );
  MUX4ND0BWP U6619 ( .I0(\vrf/regTable[4][69] ), .I1(\vrf/regTable[5][69] ), 
        .I2(\vrf/regTable[6][69] ), .I3(\vrf/regTable[7][69] ), .S0(n4939), 
        .S1(n5009), .ZN(n4435) );
  MUX2ND0BWP U6620 ( .I0(n4436), .I1(n4437), .S(n5073), .ZN(vectorData2[70])
         );
  MUX4ND0BWP U6621 ( .I0(\vrf/regTable[0][70] ), .I1(\vrf/regTable[1][70] ), 
        .I2(\vrf/regTable[2][70] ), .I3(\vrf/regTable[3][70] ), .S0(n4939), 
        .S1(n5009), .ZN(n4436) );
  MUX4ND0BWP U6622 ( .I0(\vrf/regTable[4][70] ), .I1(\vrf/regTable[5][70] ), 
        .I2(\vrf/regTable[6][70] ), .I3(\vrf/regTable[7][70] ), .S0(n4939), 
        .S1(n5009), .ZN(n4437) );
  MUX2ND0BWP U6623 ( .I0(n4438), .I1(n4439), .S(n5073), .ZN(vectorData2[71])
         );
  MUX4ND0BWP U6624 ( .I0(\vrf/regTable[0][71] ), .I1(\vrf/regTable[1][71] ), 
        .I2(\vrf/regTable[2][71] ), .I3(\vrf/regTable[3][71] ), .S0(n4939), 
        .S1(n5009), .ZN(n4438) );
  MUX4ND0BWP U6625 ( .I0(\vrf/regTable[4][71] ), .I1(\vrf/regTable[5][71] ), 
        .I2(\vrf/regTable[6][71] ), .I3(\vrf/regTable[7][71] ), .S0(n4939), 
        .S1(n5009), .ZN(n4439) );
  MUX2ND0BWP U6626 ( .I0(n4440), .I1(n4441), .S(n5069), .ZN(vectorData2[19])
         );
  MUX4ND0BWP U6627 ( .I0(\vrf/regTable[0][19] ), .I1(\vrf/regTable[1][19] ), 
        .I2(\vrf/regTable[2][19] ), .I3(\vrf/regTable[3][19] ), .S0(n4931), 
        .S1(n5001), .ZN(n4440) );
  MUX4ND0BWP U6628 ( .I0(\vrf/regTable[4][19] ), .I1(\vrf/regTable[5][19] ), 
        .I2(\vrf/regTable[6][19] ), .I3(\vrf/regTable[7][19] ), .S0(n4931), 
        .S1(n5001), .ZN(n4441) );
  MUX2ND0BWP U6629 ( .I0(n4442), .I1(n4443), .S(n5077), .ZN(vectorData2[115])
         );
  MUX4ND0BWP U6630 ( .I0(\vrf/regTable[0][115] ), .I1(\vrf/regTable[1][115] ), 
        .I2(\vrf/regTable[2][115] ), .I3(\vrf/regTable[3][115] ), .S0(n4947), 
        .S1(n5017), .ZN(n4442) );
  MUX4ND0BWP U6631 ( .I0(\vrf/regTable[4][115] ), .I1(\vrf/regTable[5][115] ), 
        .I2(\vrf/regTable[6][115] ), .I3(\vrf/regTable[7][115] ), .S0(n4947), 
        .S1(n5017), .ZN(n4443) );
  MUX2ND0BWP U6632 ( .I0(n4444), .I1(n4445), .S(n5069), .ZN(vectorData2[20])
         );
  MUX4ND0BWP U6633 ( .I0(\vrf/regTable[0][20] ), .I1(\vrf/regTable[1][20] ), 
        .I2(\vrf/regTable[2][20] ), .I3(\vrf/regTable[3][20] ), .S0(n4931), 
        .S1(n5001), .ZN(n4444) );
  MUX4ND0BWP U6634 ( .I0(\vrf/regTable[4][20] ), .I1(\vrf/regTable[5][20] ), 
        .I2(\vrf/regTable[6][20] ), .I3(\vrf/regTable[7][20] ), .S0(n4931), 
        .S1(n5001), .ZN(n4445) );
  MUX2ND0BWP U6635 ( .I0(n4446), .I1(n4447), .S(n5077), .ZN(vectorData2[116])
         );
  MUX4ND0BWP U6636 ( .I0(\vrf/regTable[0][116] ), .I1(\vrf/regTable[1][116] ), 
        .I2(\vrf/regTable[2][116] ), .I3(\vrf/regTable[3][116] ), .S0(n4947), 
        .S1(n5017), .ZN(n4446) );
  MUX4ND0BWP U6637 ( .I0(\vrf/regTable[4][116] ), .I1(\vrf/regTable[5][116] ), 
        .I2(\vrf/regTable[6][116] ), .I3(\vrf/regTable[7][116] ), .S0(n4947), 
        .S1(n5017), .ZN(n4447) );
  MUX2ND0BWP U6638 ( .I0(n4448), .I1(n4449), .S(n5080), .ZN(vectorData2[144])
         );
  MUX4ND0BWP U6639 ( .I0(\vrf/regTable[0][144] ), .I1(\vrf/regTable[1][144] ), 
        .I2(\vrf/regTable[2][144] ), .I3(\vrf/regTable[3][144] ), .S0(n4952), 
        .S1(n5022), .ZN(n4448) );
  MUX4ND0BWP U6640 ( .I0(\vrf/regTable[4][144] ), .I1(\vrf/regTable[5][144] ), 
        .I2(\vrf/regTable[6][144] ), .I3(\vrf/regTable[7][144] ), .S0(n4952), 
        .S1(n5022), .ZN(n4449) );
  MUX2ND0BWP U6641 ( .I0(n4450), .I1(n4451), .S(n5080), .ZN(vectorData2[145])
         );
  MUX4ND0BWP U6642 ( .I0(\vrf/regTable[0][145] ), .I1(\vrf/regTable[1][145] ), 
        .I2(\vrf/regTable[2][145] ), .I3(\vrf/regTable[3][145] ), .S0(n4952), 
        .S1(n5022), .ZN(n4450) );
  MUX4ND0BWP U6643 ( .I0(\vrf/regTable[4][145] ), .I1(\vrf/regTable[5][145] ), 
        .I2(\vrf/regTable[6][145] ), .I3(\vrf/regTable[7][145] ), .S0(n4952), 
        .S1(n5022), .ZN(n4451) );
  MUX2ND0BWP U6644 ( .I0(n4452), .I1(n4453), .S(n5080), .ZN(vectorData2[146])
         );
  MUX4ND0BWP U6645 ( .I0(\vrf/regTable[0][146] ), .I1(\vrf/regTable[1][146] ), 
        .I2(\vrf/regTable[2][146] ), .I3(\vrf/regTable[3][146] ), .S0(n4952), 
        .S1(n5022), .ZN(n4452) );
  MUX4ND0BWP U6646 ( .I0(\vrf/regTable[4][146] ), .I1(\vrf/regTable[5][146] ), 
        .I2(\vrf/regTable[6][146] ), .I3(\vrf/regTable[7][146] ), .S0(n4952), 
        .S1(n5022), .ZN(n4453) );
  MUX2ND0BWP U6647 ( .I0(n4454), .I1(n4455), .S(n5080), .ZN(vectorData2[149])
         );
  MUX4ND0BWP U6648 ( .I0(\vrf/regTable[0][149] ), .I1(\vrf/regTable[1][149] ), 
        .I2(\vrf/regTable[2][149] ), .I3(\vrf/regTable[3][149] ), .S0(n4952), 
        .S1(n5022), .ZN(n4454) );
  MUX4ND0BWP U6649 ( .I0(\vrf/regTable[4][149] ), .I1(\vrf/regTable[5][149] ), 
        .I2(\vrf/regTable[6][149] ), .I3(\vrf/regTable[7][149] ), .S0(n4952), 
        .S1(n5022), .ZN(n4455) );
  MUX2ND0BWP U6650 ( .I0(n4456), .I1(n4457), .S(n5080), .ZN(vectorData2[150])
         );
  MUX4ND0BWP U6651 ( .I0(\vrf/regTable[0][150] ), .I1(\vrf/regTable[1][150] ), 
        .I2(\vrf/regTable[2][150] ), .I3(\vrf/regTable[3][150] ), .S0(n4953), 
        .S1(n5023), .ZN(n4456) );
  MUX4ND0BWP U6652 ( .I0(\vrf/regTable[4][150] ), .I1(\vrf/regTable[5][150] ), 
        .I2(\vrf/regTable[6][150] ), .I3(\vrf/regTable[7][150] ), .S0(n4953), 
        .S1(n5023), .ZN(n4457) );
  MUX2ND0BWP U6653 ( .I0(n4458), .I1(n4459), .S(n5080), .ZN(vectorData2[151])
         );
  MUX4ND0BWP U6654 ( .I0(\vrf/regTable[0][151] ), .I1(\vrf/regTable[1][151] ), 
        .I2(\vrf/regTable[2][151] ), .I3(\vrf/regTable[3][151] ), .S0(n4953), 
        .S1(n5023), .ZN(n4458) );
  MUX4ND0BWP U6655 ( .I0(\vrf/regTable[4][151] ), .I1(\vrf/regTable[5][151] ), 
        .I2(\vrf/regTable[6][151] ), .I3(\vrf/regTable[7][151] ), .S0(n4953), 
        .S1(n5023), .ZN(n4459) );
  MUX2ND0BWP U6656 ( .I0(n4460), .I1(n4461), .S(n5080), .ZN(vectorData2[152])
         );
  MUX4ND0BWP U6657 ( .I0(\vrf/regTable[0][152] ), .I1(\vrf/regTable[1][152] ), 
        .I2(\vrf/regTable[2][152] ), .I3(\vrf/regTable[3][152] ), .S0(n4953), 
        .S1(n5023), .ZN(n4460) );
  MUX4ND0BWP U6658 ( .I0(\vrf/regTable[4][152] ), .I1(\vrf/regTable[5][152] ), 
        .I2(\vrf/regTable[6][152] ), .I3(\vrf/regTable[7][152] ), .S0(n4953), 
        .S1(n5023), .ZN(n4461) );
  MUX2ND0BWP U6659 ( .I0(n4462), .I1(n4463), .S(n5080), .ZN(vectorData2[153])
         );
  MUX4ND0BWP U6660 ( .I0(\vrf/regTable[0][153] ), .I1(\vrf/regTable[1][153] ), 
        .I2(\vrf/regTable[2][153] ), .I3(\vrf/regTable[3][153] ), .S0(n4953), 
        .S1(n5023), .ZN(n4462) );
  MUX4ND0BWP U6661 ( .I0(\vrf/regTable[4][153] ), .I1(\vrf/regTable[5][153] ), 
        .I2(\vrf/regTable[6][153] ), .I3(\vrf/regTable[7][153] ), .S0(n4953), 
        .S1(n5023), .ZN(n4463) );
  MUX2ND0BWP U6662 ( .I0(n4464), .I1(n4465), .S(n5080), .ZN(vectorData2[154])
         );
  MUX4ND0BWP U6663 ( .I0(\vrf/regTable[0][154] ), .I1(\vrf/regTable[1][154] ), 
        .I2(\vrf/regTable[2][154] ), .I3(\vrf/regTable[3][154] ), .S0(n4953), 
        .S1(n5023), .ZN(n4464) );
  MUX4ND0BWP U6664 ( .I0(\vrf/regTable[4][154] ), .I1(\vrf/regTable[5][154] ), 
        .I2(\vrf/regTable[6][154] ), .I3(\vrf/regTable[7][154] ), .S0(n4953), 
        .S1(n5023), .ZN(n4465) );
  MUX2ND0BWP U6665 ( .I0(n4466), .I1(n4467), .S(n5080), .ZN(vectorData2[155])
         );
  MUX4ND0BWP U6666 ( .I0(\vrf/regTable[0][155] ), .I1(\vrf/regTable[1][155] ), 
        .I2(\vrf/regTable[2][155] ), .I3(\vrf/regTable[3][155] ), .S0(n4953), 
        .S1(n5023), .ZN(n4466) );
  MUX4ND0BWP U6667 ( .I0(\vrf/regTable[4][155] ), .I1(\vrf/regTable[5][155] ), 
        .I2(\vrf/regTable[6][155] ), .I3(\vrf/regTable[7][155] ), .S0(n4953), 
        .S1(n5023), .ZN(n4467) );
  MUX2ND0BWP U6668 ( .I0(n4468), .I1(n4469), .S(n5081), .ZN(vectorData2[156])
         );
  MUX4ND0BWP U6669 ( .I0(\vrf/regTable[0][156] ), .I1(\vrf/regTable[1][156] ), 
        .I2(\vrf/regTable[2][156] ), .I3(\vrf/regTable[3][156] ), .S0(n4954), 
        .S1(n5024), .ZN(n4468) );
  MUX4ND0BWP U6670 ( .I0(\vrf/regTable[4][156] ), .I1(\vrf/regTable[5][156] ), 
        .I2(\vrf/regTable[6][156] ), .I3(\vrf/regTable[7][156] ), .S0(n4954), 
        .S1(n5024), .ZN(n4469) );
  MUX2ND0BWP U6671 ( .I0(n4470), .I1(n4471), .S(n5081), .ZN(vectorData2[157])
         );
  MUX4ND0BWP U6672 ( .I0(\vrf/regTable[0][157] ), .I1(\vrf/regTable[1][157] ), 
        .I2(\vrf/regTable[2][157] ), .I3(\vrf/regTable[3][157] ), .S0(n4954), 
        .S1(n5024), .ZN(n4470) );
  MUX4ND0BWP U6673 ( .I0(\vrf/regTable[4][157] ), .I1(\vrf/regTable[5][157] ), 
        .I2(\vrf/regTable[6][157] ), .I3(\vrf/regTable[7][157] ), .S0(n4954), 
        .S1(n5024), .ZN(n4471) );
  MUX2ND0BWP U6674 ( .I0(n4472), .I1(n4473), .S(n5081), .ZN(vectorData2[158])
         );
  MUX4ND0BWP U6675 ( .I0(\vrf/regTable[0][158] ), .I1(\vrf/regTable[1][158] ), 
        .I2(\vrf/regTable[2][158] ), .I3(\vrf/regTable[3][158] ), .S0(n4954), 
        .S1(n5024), .ZN(n4472) );
  MUX4ND0BWP U6676 ( .I0(\vrf/regTable[4][158] ), .I1(\vrf/regTable[5][158] ), 
        .I2(\vrf/regTable[6][158] ), .I3(\vrf/regTable[7][158] ), .S0(n4954), 
        .S1(n5024), .ZN(n4473) );
  MUX2ND0BWP U6677 ( .I0(n4474), .I1(n4475), .S(n5081), .ZN(vectorData2[159])
         );
  MUX4ND0BWP U6678 ( .I0(\vrf/regTable[0][159] ), .I1(\vrf/regTable[1][159] ), 
        .I2(\vrf/regTable[2][159] ), .I3(\vrf/regTable[3][159] ), .S0(n4954), 
        .S1(n5024), .ZN(n4474) );
  MUX4ND0BWP U6679 ( .I0(\vrf/regTable[4][159] ), .I1(\vrf/regTable[5][159] ), 
        .I2(\vrf/regTable[6][159] ), .I3(\vrf/regTable[7][159] ), .S0(n4954), 
        .S1(n5024), .ZN(n4475) );
  MUX2ND0BWP U6680 ( .I0(n4476), .I1(n4477), .S(n5084), .ZN(vectorData2[192])
         );
  MUX4ND0BWP U6681 ( .I0(\vrf/regTable[0][192] ), .I1(\vrf/regTable[1][192] ), 
        .I2(\vrf/regTable[2][192] ), .I3(\vrf/regTable[3][192] ), .S0(n4960), 
        .S1(n5030), .ZN(n4476) );
  MUX4ND0BWP U6682 ( .I0(\vrf/regTable[4][192] ), .I1(\vrf/regTable[5][192] ), 
        .I2(\vrf/regTable[6][192] ), .I3(\vrf/regTable[7][192] ), .S0(n4960), 
        .S1(n5030), .ZN(n4477) );
  MUX2ND0BWP U6683 ( .I0(n4478), .I1(n4479), .S(n5070), .ZN(vectorData2[32])
         );
  MUX4ND0BWP U6684 ( .I0(\vrf/regTable[0][32] ), .I1(\vrf/regTable[1][32] ), 
        .I2(\vrf/regTable[2][32] ), .I3(\vrf/regTable[3][32] ), .S0(n4933), 
        .S1(n5003), .ZN(n4478) );
  MUX4ND0BWP U6685 ( .I0(\vrf/regTable[4][32] ), .I1(\vrf/regTable[5][32] ), 
        .I2(\vrf/regTable[6][32] ), .I3(\vrf/regTable[7][32] ), .S0(n4933), 
        .S1(n5003), .ZN(n4479) );
  MUX2ND0BWP U6686 ( .I0(n4480), .I1(n4481), .S(n5084), .ZN(vectorData2[193])
         );
  MUX4ND0BWP U6687 ( .I0(\vrf/regTable[0][193] ), .I1(\vrf/regTable[1][193] ), 
        .I2(\vrf/regTable[2][193] ), .I3(\vrf/regTable[3][193] ), .S0(n4960), 
        .S1(n5030), .ZN(n4480) );
  MUX4ND0BWP U6688 ( .I0(\vrf/regTable[4][193] ), .I1(\vrf/regTable[5][193] ), 
        .I2(\vrf/regTable[6][193] ), .I3(\vrf/regTable[7][193] ), .S0(n4960), 
        .S1(n5030), .ZN(n4481) );
  MUX2ND0BWP U6689 ( .I0(n4482), .I1(n4483), .S(n5070), .ZN(vectorData2[33])
         );
  MUX4ND0BWP U6690 ( .I0(\vrf/regTable[0][33] ), .I1(\vrf/regTable[1][33] ), 
        .I2(\vrf/regTable[2][33] ), .I3(\vrf/regTable[3][33] ), .S0(n4933), 
        .S1(n5003), .ZN(n4482) );
  MUX4ND0BWP U6691 ( .I0(\vrf/regTable[4][33] ), .I1(\vrf/regTable[5][33] ), 
        .I2(\vrf/regTable[6][33] ), .I3(\vrf/regTable[7][33] ), .S0(n4933), 
        .S1(n5003), .ZN(n4483) );
  MUX2ND0BWP U6692 ( .I0(n4484), .I1(n4485), .S(n5084), .ZN(vectorData2[200])
         );
  MUX4ND0BWP U6693 ( .I0(\vrf/regTable[0][200] ), .I1(\vrf/regTable[1][200] ), 
        .I2(\vrf/regTable[2][200] ), .I3(\vrf/regTable[3][200] ), .S0(n4961), 
        .S1(n5031), .ZN(n4484) );
  MUX4ND0BWP U6694 ( .I0(\vrf/regTable[4][200] ), .I1(\vrf/regTable[5][200] ), 
        .I2(\vrf/regTable[6][200] ), .I3(\vrf/regTable[7][200] ), .S0(n4961), 
        .S1(n5031), .ZN(n4485) );
  MUX2ND0BWP U6695 ( .I0(n4486), .I1(n4487), .S(n5071), .ZN(vectorData2[40])
         );
  MUX4ND0BWP U6696 ( .I0(\vrf/regTable[0][40] ), .I1(\vrf/regTable[1][40] ), 
        .I2(\vrf/regTable[2][40] ), .I3(\vrf/regTable[3][40] ), .S0(n4934), 
        .S1(n5004), .ZN(n4486) );
  MUX4ND0BWP U6697 ( .I0(\vrf/regTable[4][40] ), .I1(\vrf/regTable[5][40] ), 
        .I2(\vrf/regTable[6][40] ), .I3(\vrf/regTable[7][40] ), .S0(n4934), 
        .S1(n5004), .ZN(n4487) );
  MUX2ND0BWP U6698 ( .I0(n4488), .I1(n4489), .S(n5084), .ZN(vectorData2[201])
         );
  MUX4ND0BWP U6699 ( .I0(\vrf/regTable[0][201] ), .I1(\vrf/regTable[1][201] ), 
        .I2(\vrf/regTable[2][201] ), .I3(\vrf/regTable[3][201] ), .S0(n4961), 
        .S1(n5031), .ZN(n4488) );
  MUX4ND0BWP U6700 ( .I0(\vrf/regTable[4][201] ), .I1(\vrf/regTable[5][201] ), 
        .I2(\vrf/regTable[6][201] ), .I3(\vrf/regTable[7][201] ), .S0(n4961), 
        .S1(n5031), .ZN(n4489) );
  MUX2ND0BWP U6701 ( .I0(n4490), .I1(n4491), .S(n5071), .ZN(vectorData2[41])
         );
  MUX4ND0BWP U6702 ( .I0(\vrf/regTable[0][41] ), .I1(\vrf/regTable[1][41] ), 
        .I2(\vrf/regTable[2][41] ), .I3(\vrf/regTable[3][41] ), .S0(n4934), 
        .S1(n5004), .ZN(n4490) );
  MUX4ND0BWP U6703 ( .I0(\vrf/regTable[4][41] ), .I1(\vrf/regTable[5][41] ), 
        .I2(\vrf/regTable[6][41] ), .I3(\vrf/regTable[7][41] ), .S0(n4934), 
        .S1(n5004), .ZN(n4491) );
  MUX2ND0BWP U6704 ( .I0(n4492), .I1(n4493), .S(n5084), .ZN(vectorData2[202])
         );
  MUX4ND0BWP U6705 ( .I0(\vrf/regTable[0][202] ), .I1(\vrf/regTable[1][202] ), 
        .I2(\vrf/regTable[2][202] ), .I3(\vrf/regTable[3][202] ), .S0(n4961), 
        .S1(n5031), .ZN(n4492) );
  MUX4ND0BWP U6706 ( .I0(\vrf/regTable[4][202] ), .I1(\vrf/regTable[5][202] ), 
        .I2(\vrf/regTable[6][202] ), .I3(\vrf/regTable[7][202] ), .S0(n4961), 
        .S1(n5031), .ZN(n4493) );
  MUX2ND0BWP U6707 ( .I0(n4494), .I1(n4495), .S(n5071), .ZN(vectorData2[42])
         );
  MUX4ND0BWP U6708 ( .I0(\vrf/regTable[0][42] ), .I1(\vrf/regTable[1][42] ), 
        .I2(\vrf/regTable[2][42] ), .I3(\vrf/regTable[3][42] ), .S0(n4935), 
        .S1(n5005), .ZN(n4494) );
  MUX4ND0BWP U6709 ( .I0(\vrf/regTable[4][42] ), .I1(\vrf/regTable[5][42] ), 
        .I2(\vrf/regTable[6][42] ), .I3(\vrf/regTable[7][42] ), .S0(n4935), 
        .S1(n5005), .ZN(n4495) );
  MUX2ND0BWP U6710 ( .I0(n4496), .I1(n4497), .S(n5084), .ZN(vectorData2[203])
         );
  MUX4ND0BWP U6711 ( .I0(\vrf/regTable[0][203] ), .I1(\vrf/regTable[1][203] ), 
        .I2(\vrf/regTable[2][203] ), .I3(\vrf/regTable[3][203] ), .S0(n4961), 
        .S1(n5031), .ZN(n4496) );
  MUX4ND0BWP U6712 ( .I0(\vrf/regTable[4][203] ), .I1(\vrf/regTable[5][203] ), 
        .I2(\vrf/regTable[6][203] ), .I3(\vrf/regTable[7][203] ), .S0(n4961), 
        .S1(n5031), .ZN(n4497) );
  MUX2ND0BWP U6713 ( .I0(n4498), .I1(n4499), .S(n5071), .ZN(vectorData2[43])
         );
  MUX4ND0BWP U6714 ( .I0(\vrf/regTable[0][43] ), .I1(\vrf/regTable[1][43] ), 
        .I2(\vrf/regTable[2][43] ), .I3(\vrf/regTable[3][43] ), .S0(n4935), 
        .S1(n5005), .ZN(n4498) );
  MUX4ND0BWP U6715 ( .I0(\vrf/regTable[4][43] ), .I1(\vrf/regTable[5][43] ), 
        .I2(\vrf/regTable[6][43] ), .I3(\vrf/regTable[7][43] ), .S0(n4935), 
        .S1(n5005), .ZN(n4499) );
  MUX2ND0BWP U6716 ( .I0(n4500), .I1(n4501), .S(n5085), .ZN(vectorData2[204])
         );
  MUX4ND0BWP U6717 ( .I0(\vrf/regTable[0][204] ), .I1(\vrf/regTable[1][204] ), 
        .I2(\vrf/regTable[2][204] ), .I3(\vrf/regTable[3][204] ), .S0(n4962), 
        .S1(n5032), .ZN(n4500) );
  MUX4ND0BWP U6718 ( .I0(\vrf/regTable[4][204] ), .I1(\vrf/regTable[5][204] ), 
        .I2(\vrf/regTable[6][204] ), .I3(\vrf/regTable[7][204] ), .S0(n4962), 
        .S1(n5032), .ZN(n4501) );
  MUX2ND0BWP U6719 ( .I0(n4502), .I1(n4503), .S(n5071), .ZN(vectorData2[44])
         );
  MUX4ND0BWP U6720 ( .I0(\vrf/regTable[0][44] ), .I1(\vrf/regTable[1][44] ), 
        .I2(\vrf/regTable[2][44] ), .I3(\vrf/regTable[3][44] ), .S0(n4935), 
        .S1(n5005), .ZN(n4502) );
  MUX4ND0BWP U6721 ( .I0(\vrf/regTable[4][44] ), .I1(\vrf/regTable[5][44] ), 
        .I2(\vrf/regTable[6][44] ), .I3(\vrf/regTable[7][44] ), .S0(n4935), 
        .S1(n5005), .ZN(n4503) );
  MUX2ND0BWP U6722 ( .I0(n4504), .I1(n4505), .S(n5085), .ZN(vectorData2[205])
         );
  MUX4ND0BWP U6723 ( .I0(\vrf/regTable[0][205] ), .I1(\vrf/regTable[1][205] ), 
        .I2(\vrf/regTable[2][205] ), .I3(\vrf/regTable[3][205] ), .S0(n4962), 
        .S1(n5032), .ZN(n4504) );
  MUX4ND0BWP U6724 ( .I0(\vrf/regTable[4][205] ), .I1(\vrf/regTable[5][205] ), 
        .I2(\vrf/regTable[6][205] ), .I3(\vrf/regTable[7][205] ), .S0(n4962), 
        .S1(n5032), .ZN(n4505) );
  MUX2ND0BWP U6725 ( .I0(n4506), .I1(n4507), .S(n5071), .ZN(vectorData2[45])
         );
  MUX4ND0BWP U6726 ( .I0(\vrf/regTable[0][45] ), .I1(\vrf/regTable[1][45] ), 
        .I2(\vrf/regTable[2][45] ), .I3(\vrf/regTable[3][45] ), .S0(n4935), 
        .S1(n5005), .ZN(n4506) );
  MUX4ND0BWP U6727 ( .I0(\vrf/regTable[4][45] ), .I1(\vrf/regTable[5][45] ), 
        .I2(\vrf/regTable[6][45] ), .I3(\vrf/regTable[7][45] ), .S0(n4935), 
        .S1(n5005), .ZN(n4507) );
  MUX2ND0BWP U6728 ( .I0(n4508), .I1(n4509), .S(n5085), .ZN(vectorData2[206])
         );
  MUX4ND0BWP U6729 ( .I0(\vrf/regTable[0][206] ), .I1(\vrf/regTable[1][206] ), 
        .I2(\vrf/regTable[2][206] ), .I3(\vrf/regTable[3][206] ), .S0(n4962), 
        .S1(n5032), .ZN(n4508) );
  MUX4ND0BWP U6730 ( .I0(\vrf/regTable[4][206] ), .I1(\vrf/regTable[5][206] ), 
        .I2(\vrf/regTable[6][206] ), .I3(\vrf/regTable[7][206] ), .S0(n4962), 
        .S1(n5032), .ZN(n4509) );
  MUX2ND0BWP U6731 ( .I0(n4510), .I1(n4511), .S(n5071), .ZN(vectorData2[46])
         );
  MUX4ND0BWP U6732 ( .I0(\vrf/regTable[0][46] ), .I1(\vrf/regTable[1][46] ), 
        .I2(\vrf/regTable[2][46] ), .I3(\vrf/regTable[3][46] ), .S0(n4935), 
        .S1(n5005), .ZN(n4510) );
  MUX4ND0BWP U6733 ( .I0(\vrf/regTable[4][46] ), .I1(\vrf/regTable[5][46] ), 
        .I2(\vrf/regTable[6][46] ), .I3(\vrf/regTable[7][46] ), .S0(n4935), 
        .S1(n5005), .ZN(n4511) );
  MUX2ND0BWP U6734 ( .I0(n4512), .I1(n4513), .S(n5085), .ZN(vectorData2[207])
         );
  MUX4ND0BWP U6735 ( .I0(\vrf/regTable[0][207] ), .I1(\vrf/regTable[1][207] ), 
        .I2(\vrf/regTable[2][207] ), .I3(\vrf/regTable[3][207] ), .S0(n4962), 
        .S1(n5032), .ZN(n4512) );
  MUX4ND0BWP U6736 ( .I0(\vrf/regTable[4][207] ), .I1(\vrf/regTable[5][207] ), 
        .I2(\vrf/regTable[6][207] ), .I3(\vrf/regTable[7][207] ), .S0(n4962), 
        .S1(n5032), .ZN(n4513) );
  MUX2ND0BWP U6737 ( .I0(n4514), .I1(n4515), .S(n5071), .ZN(vectorData2[47])
         );
  MUX4ND0BWP U6738 ( .I0(\vrf/regTable[0][47] ), .I1(\vrf/regTable[1][47] ), 
        .I2(\vrf/regTable[2][47] ), .I3(\vrf/regTable[3][47] ), .S0(n4935), 
        .S1(n5005), .ZN(n4514) );
  MUX4ND0BWP U6739 ( .I0(\vrf/regTable[4][47] ), .I1(\vrf/regTable[5][47] ), 
        .I2(\vrf/regTable[6][47] ), .I3(\vrf/regTable[7][47] ), .S0(n4935), 
        .S1(n5005), .ZN(n4515) );
  MUX2ND0BWP U6740 ( .I0(n4516), .I1(n4517), .S(n5084), .ZN(vectorData2[194])
         );
  MUX4ND0BWP U6741 ( .I0(\vrf/regTable[0][194] ), .I1(\vrf/regTable[1][194] ), 
        .I2(\vrf/regTable[2][194] ), .I3(\vrf/regTable[3][194] ), .S0(n4960), 
        .S1(n5030), .ZN(n4516) );
  MUX4ND0BWP U6742 ( .I0(\vrf/regTable[4][194] ), .I1(\vrf/regTable[5][194] ), 
        .I2(\vrf/regTable[6][194] ), .I3(\vrf/regTable[7][194] ), .S0(n4960), 
        .S1(n5030), .ZN(n4517) );
  MUX2ND0BWP U6743 ( .I0(n4518), .I1(n4519), .S(n5070), .ZN(vectorData2[34])
         );
  MUX4ND0BWP U6744 ( .I0(\vrf/regTable[0][34] ), .I1(\vrf/regTable[1][34] ), 
        .I2(\vrf/regTable[2][34] ), .I3(\vrf/regTable[3][34] ), .S0(n4933), 
        .S1(n5003), .ZN(n4518) );
  MUX4ND0BWP U6745 ( .I0(\vrf/regTable[4][34] ), .I1(\vrf/regTable[5][34] ), 
        .I2(\vrf/regTable[6][34] ), .I3(\vrf/regTable[7][34] ), .S0(n4933), 
        .S1(n5003), .ZN(n4519) );
  MUX2ND0BWP U6746 ( .I0(n4520), .I1(n4521), .S(n5084), .ZN(vectorData2[197])
         );
  MUX4ND0BWP U6747 ( .I0(\vrf/regTable[0][197] ), .I1(\vrf/regTable[1][197] ), 
        .I2(\vrf/regTable[2][197] ), .I3(\vrf/regTable[3][197] ), .S0(n4960), 
        .S1(n5030), .ZN(n4520) );
  MUX4ND0BWP U6748 ( .I0(\vrf/regTable[4][197] ), .I1(\vrf/regTable[5][197] ), 
        .I2(\vrf/regTable[6][197] ), .I3(\vrf/regTable[7][197] ), .S0(n4960), 
        .S1(n5030), .ZN(n4521) );
  MUX2ND0BWP U6749 ( .I0(n4522), .I1(n4523), .S(n5071), .ZN(vectorData2[37])
         );
  MUX4ND0BWP U6750 ( .I0(\vrf/regTable[0][37] ), .I1(\vrf/regTable[1][37] ), 
        .I2(\vrf/regTable[2][37] ), .I3(\vrf/regTable[3][37] ), .S0(n4934), 
        .S1(n5004), .ZN(n4522) );
  MUX4ND0BWP U6751 ( .I0(\vrf/regTable[4][37] ), .I1(\vrf/regTable[5][37] ), 
        .I2(\vrf/regTable[6][37] ), .I3(\vrf/regTable[7][37] ), .S0(n4934), 
        .S1(n5004), .ZN(n4523) );
  MUX2ND0BWP U6752 ( .I0(n4524), .I1(n4525), .S(n5084), .ZN(vectorData2[198])
         );
  MUX4ND0BWP U6753 ( .I0(\vrf/regTable[0][198] ), .I1(\vrf/regTable[1][198] ), 
        .I2(\vrf/regTable[2][198] ), .I3(\vrf/regTable[3][198] ), .S0(n4961), 
        .S1(n5031), .ZN(n4524) );
  MUX4ND0BWP U6754 ( .I0(\vrf/regTable[4][198] ), .I1(\vrf/regTable[5][198] ), 
        .I2(\vrf/regTable[6][198] ), .I3(\vrf/regTable[7][198] ), .S0(n4961), 
        .S1(n5031), .ZN(n4525) );
  MUX2ND0BWP U6755 ( .I0(n4526), .I1(n4527), .S(n5071), .ZN(vectorData2[38])
         );
  MUX4ND0BWP U6756 ( .I0(\vrf/regTable[0][38] ), .I1(\vrf/regTable[1][38] ), 
        .I2(\vrf/regTable[2][38] ), .I3(\vrf/regTable[3][38] ), .S0(n4934), 
        .S1(n5004), .ZN(n4526) );
  MUX4ND0BWP U6757 ( .I0(\vrf/regTable[4][38] ), .I1(\vrf/regTable[5][38] ), 
        .I2(\vrf/regTable[6][38] ), .I3(\vrf/regTable[7][38] ), .S0(n4934), 
        .S1(n5004), .ZN(n4527) );
  MUX2ND0BWP U6758 ( .I0(n4528), .I1(n4529), .S(n5084), .ZN(vectorData2[199])
         );
  MUX4ND0BWP U6759 ( .I0(\vrf/regTable[0][199] ), .I1(\vrf/regTable[1][199] ), 
        .I2(\vrf/regTable[2][199] ), .I3(\vrf/regTable[3][199] ), .S0(n4961), 
        .S1(n5031), .ZN(n4528) );
  MUX4ND0BWP U6760 ( .I0(\vrf/regTable[4][199] ), .I1(\vrf/regTable[5][199] ), 
        .I2(\vrf/regTable[6][199] ), .I3(\vrf/regTable[7][199] ), .S0(n4961), 
        .S1(n5031), .ZN(n4529) );
  MUX2ND0BWP U6761 ( .I0(n4530), .I1(n4531), .S(n5071), .ZN(vectorData2[39])
         );
  MUX4ND0BWP U6762 ( .I0(\vrf/regTable[0][39] ), .I1(\vrf/regTable[1][39] ), 
        .I2(\vrf/regTable[2][39] ), .I3(\vrf/regTable[3][39] ), .S0(n4934), 
        .S1(n5004), .ZN(n4530) );
  MUX4ND0BWP U6763 ( .I0(\vrf/regTable[4][39] ), .I1(\vrf/regTable[5][39] ), 
        .I2(\vrf/regTable[6][39] ), .I3(\vrf/regTable[7][39] ), .S0(n4934), 
        .S1(n5004), .ZN(n4531) );
  MUX2ND0BWP U6764 ( .I0(n4532), .I1(n4533), .S(n5080), .ZN(vectorData2[147])
         );
  MUX4ND0BWP U6765 ( .I0(\vrf/regTable[0][147] ), .I1(\vrf/regTable[1][147] ), 
        .I2(\vrf/regTable[2][147] ), .I3(\vrf/regTable[3][147] ), .S0(n4952), 
        .S1(n5022), .ZN(n4532) );
  MUX4ND0BWP U6766 ( .I0(\vrf/regTable[4][147] ), .I1(\vrf/regTable[5][147] ), 
        .I2(\vrf/regTable[6][147] ), .I3(\vrf/regTable[7][147] ), .S0(n4952), 
        .S1(n5022), .ZN(n4533) );
  MUX2ND0BWP U6767 ( .I0(n4534), .I1(n4535), .S(n5080), .ZN(vectorData2[148])
         );
  MUX4ND0BWP U6768 ( .I0(\vrf/regTable[0][148] ), .I1(\vrf/regTable[1][148] ), 
        .I2(\vrf/regTable[2][148] ), .I3(\vrf/regTable[3][148] ), .S0(n4952), 
        .S1(n5022), .ZN(n4534) );
  MUX4ND0BWP U6769 ( .I0(\vrf/regTable[4][148] ), .I1(\vrf/regTable[5][148] ), 
        .I2(\vrf/regTable[6][148] ), .I3(\vrf/regTable[7][148] ), .S0(n4952), 
        .S1(n5022), .ZN(n4535) );
  MUX2ND0BWP U6770 ( .I0(n4536), .I1(n4537), .S(n5076), .ZN(vectorData2[96])
         );
  MUX4ND0BWP U6771 ( .I0(\vrf/regTable[0][96] ), .I1(\vrf/regTable[1][96] ), 
        .I2(\vrf/regTable[2][96] ), .I3(\vrf/regTable[3][96] ), .S0(n4944), 
        .S1(n5014), .ZN(n4536) );
  MUX4ND0BWP U6772 ( .I0(\vrf/regTable[4][96] ), .I1(\vrf/regTable[5][96] ), 
        .I2(\vrf/regTable[6][96] ), .I3(\vrf/regTable[7][96] ), .S0(n4944), 
        .S1(n5014), .ZN(n4537) );
  MUX2ND0BWP U6773 ( .I0(n4538), .I1(n4539), .S(n5076), .ZN(vectorData2[97])
         );
  MUX4ND0BWP U6774 ( .I0(\vrf/regTable[0][97] ), .I1(\vrf/regTable[1][97] ), 
        .I2(\vrf/regTable[2][97] ), .I3(\vrf/regTable[3][97] ), .S0(n4944), 
        .S1(n5014), .ZN(n4538) );
  MUX4ND0BWP U6775 ( .I0(\vrf/regTable[4][97] ), .I1(\vrf/regTable[5][97] ), 
        .I2(\vrf/regTable[6][97] ), .I3(\vrf/regTable[7][97] ), .S0(n4944), 
        .S1(n5014), .ZN(n4539) );
  MUX2ND0BWP U6776 ( .I0(n4540), .I1(n4541), .S(n5076), .ZN(vectorData2[104])
         );
  MUX4ND0BWP U6777 ( .I0(\vrf/regTable[0][104] ), .I1(\vrf/regTable[1][104] ), 
        .I2(\vrf/regTable[2][104] ), .I3(\vrf/regTable[3][104] ), .S0(n4945), 
        .S1(n5015), .ZN(n4540) );
  MUX4ND0BWP U6778 ( .I0(\vrf/regTable[4][104] ), .I1(\vrf/regTable[5][104] ), 
        .I2(\vrf/regTable[6][104] ), .I3(\vrf/regTable[7][104] ), .S0(n4945), 
        .S1(n5015), .ZN(n4541) );
  MUX2ND0BWP U6779 ( .I0(n4542), .I1(n4543), .S(n5076), .ZN(vectorData2[105])
         );
  MUX4ND0BWP U6780 ( .I0(\vrf/regTable[0][105] ), .I1(\vrf/regTable[1][105] ), 
        .I2(\vrf/regTable[2][105] ), .I3(\vrf/regTable[3][105] ), .S0(n4945), 
        .S1(n5015), .ZN(n4542) );
  MUX4ND0BWP U6781 ( .I0(\vrf/regTable[4][105] ), .I1(\vrf/regTable[5][105] ), 
        .I2(\vrf/regTable[6][105] ), .I3(\vrf/regTable[7][105] ), .S0(n4945), 
        .S1(n5015), .ZN(n4543) );
  MUX2ND0BWP U6782 ( .I0(n4544), .I1(n4545), .S(n5076), .ZN(vectorData2[106])
         );
  MUX4ND0BWP U6783 ( .I0(\vrf/regTable[0][106] ), .I1(\vrf/regTable[1][106] ), 
        .I2(\vrf/regTable[2][106] ), .I3(\vrf/regTable[3][106] ), .S0(n4945), 
        .S1(n5015), .ZN(n4544) );
  MUX4ND0BWP U6784 ( .I0(\vrf/regTable[4][106] ), .I1(\vrf/regTable[5][106] ), 
        .I2(\vrf/regTable[6][106] ), .I3(\vrf/regTable[7][106] ), .S0(n4945), 
        .S1(n5015), .ZN(n4545) );
  MUX2ND0BWP U6785 ( .I0(n4546), .I1(n4547), .S(n5076), .ZN(vectorData2[107])
         );
  MUX4ND0BWP U6786 ( .I0(\vrf/regTable[0][107] ), .I1(\vrf/regTable[1][107] ), 
        .I2(\vrf/regTable[2][107] ), .I3(\vrf/regTable[3][107] ), .S0(n4945), 
        .S1(n5015), .ZN(n4546) );
  MUX4ND0BWP U6787 ( .I0(\vrf/regTable[4][107] ), .I1(\vrf/regTable[5][107] ), 
        .I2(\vrf/regTable[6][107] ), .I3(\vrf/regTable[7][107] ), .S0(n4945), 
        .S1(n5015), .ZN(n4547) );
  MUX2ND0BWP U6788 ( .I0(n4548), .I1(n4549), .S(n5077), .ZN(vectorData2[108])
         );
  MUX4ND0BWP U6789 ( .I0(\vrf/regTable[0][108] ), .I1(\vrf/regTable[1][108] ), 
        .I2(\vrf/regTable[2][108] ), .I3(\vrf/regTable[3][108] ), .S0(n4946), 
        .S1(n5016), .ZN(n4548) );
  MUX4ND0BWP U6790 ( .I0(\vrf/regTable[4][108] ), .I1(\vrf/regTable[5][108] ), 
        .I2(\vrf/regTable[6][108] ), .I3(\vrf/regTable[7][108] ), .S0(n4946), 
        .S1(n5016), .ZN(n4549) );
  MUX2ND0BWP U6791 ( .I0(n4550), .I1(n4551), .S(n5077), .ZN(vectorData2[109])
         );
  MUX4ND0BWP U6792 ( .I0(\vrf/regTable[0][109] ), .I1(\vrf/regTable[1][109] ), 
        .I2(\vrf/regTable[2][109] ), .I3(\vrf/regTable[3][109] ), .S0(n4946), 
        .S1(n5016), .ZN(n4550) );
  MUX4ND0BWP U6793 ( .I0(\vrf/regTable[4][109] ), .I1(\vrf/regTable[5][109] ), 
        .I2(\vrf/regTable[6][109] ), .I3(\vrf/regTable[7][109] ), .S0(n4946), 
        .S1(n5016), .ZN(n4551) );
  MUX2ND0BWP U6794 ( .I0(n4552), .I1(n4553), .S(n5077), .ZN(vectorData2[110])
         );
  MUX4ND0BWP U6795 ( .I0(\vrf/regTable[0][110] ), .I1(\vrf/regTable[1][110] ), 
        .I2(\vrf/regTable[2][110] ), .I3(\vrf/regTable[3][110] ), .S0(n4946), 
        .S1(n5016), .ZN(n4552) );
  MUX4ND0BWP U6796 ( .I0(\vrf/regTable[4][110] ), .I1(\vrf/regTable[5][110] ), 
        .I2(\vrf/regTable[6][110] ), .I3(\vrf/regTable[7][110] ), .S0(n4946), 
        .S1(n5016), .ZN(n4553) );
  MUX2ND0BWP U6797 ( .I0(n4554), .I1(n4555), .S(n5077), .ZN(vectorData2[111])
         );
  MUX4ND0BWP U6798 ( .I0(\vrf/regTable[0][111] ), .I1(\vrf/regTable[1][111] ), 
        .I2(\vrf/regTable[2][111] ), .I3(\vrf/regTable[3][111] ), .S0(n4946), 
        .S1(n5016), .ZN(n4554) );
  MUX4ND0BWP U6799 ( .I0(\vrf/regTable[4][111] ), .I1(\vrf/regTable[5][111] ), 
        .I2(\vrf/regTable[6][111] ), .I3(\vrf/regTable[7][111] ), .S0(n4946), 
        .S1(n5016), .ZN(n4555) );
  MUX2ND0BWP U6800 ( .I0(n4556), .I1(n4557), .S(n5076), .ZN(vectorData2[98])
         );
  MUX4ND0BWP U6801 ( .I0(\vrf/regTable[0][98] ), .I1(\vrf/regTable[1][98] ), 
        .I2(\vrf/regTable[2][98] ), .I3(\vrf/regTable[3][98] ), .S0(n4944), 
        .S1(n5014), .ZN(n4556) );
  MUX4ND0BWP U6802 ( .I0(\vrf/regTable[4][98] ), .I1(\vrf/regTable[5][98] ), 
        .I2(\vrf/regTable[6][98] ), .I3(\vrf/regTable[7][98] ), .S0(n4944), 
        .S1(n5014), .ZN(n4557) );
  MUX2ND0BWP U6803 ( .I0(n4558), .I1(n4559), .S(n5076), .ZN(vectorData2[101])
         );
  MUX4ND0BWP U6804 ( .I0(\vrf/regTable[0][101] ), .I1(\vrf/regTable[1][101] ), 
        .I2(\vrf/regTable[2][101] ), .I3(\vrf/regTable[3][101] ), .S0(n4944), 
        .S1(n5014), .ZN(n4558) );
  MUX4ND0BWP U6805 ( .I0(\vrf/regTable[4][101] ), .I1(\vrf/regTable[5][101] ), 
        .I2(\vrf/regTable[6][101] ), .I3(\vrf/regTable[7][101] ), .S0(n4944), 
        .S1(n5014), .ZN(n4559) );
  MUX2ND0BWP U6806 ( .I0(n4560), .I1(n4561), .S(n5076), .ZN(vectorData2[102])
         );
  MUX4ND0BWP U6807 ( .I0(\vrf/regTable[0][102] ), .I1(\vrf/regTable[1][102] ), 
        .I2(\vrf/regTable[2][102] ), .I3(\vrf/regTable[3][102] ), .S0(n4945), 
        .S1(n5015), .ZN(n4560) );
  MUX4ND0BWP U6808 ( .I0(\vrf/regTable[4][102] ), .I1(\vrf/regTable[5][102] ), 
        .I2(\vrf/regTable[6][102] ), .I3(\vrf/regTable[7][102] ), .S0(n4945), 
        .S1(n5015), .ZN(n4561) );
  MUX2ND0BWP U6809 ( .I0(n4562), .I1(n4563), .S(n5076), .ZN(vectorData2[103])
         );
  MUX4ND0BWP U6810 ( .I0(\vrf/regTable[0][103] ), .I1(\vrf/regTable[1][103] ), 
        .I2(\vrf/regTable[2][103] ), .I3(\vrf/regTable[3][103] ), .S0(n4945), 
        .S1(n5015), .ZN(n4562) );
  MUX4ND0BWP U6811 ( .I0(\vrf/regTable[4][103] ), .I1(\vrf/regTable[5][103] ), 
        .I2(\vrf/regTable[6][103] ), .I3(\vrf/regTable[7][103] ), .S0(n4945), 
        .S1(n5015), .ZN(n4563) );
  MUX2ND0BWP U6812 ( .I0(n4564), .I1(n4565), .S(n4914), .ZN(scalarData1[0]) );
  MUX4ND0BWP U6813 ( .I0(\srf/regTable[0][0] ), .I1(\srf/regTable[1][0] ), 
        .I2(\srf/regTable[2][0] ), .I3(\srf/regTable[3][0] ), .S0(n4795), .S1(
        n4865), .ZN(n4564) );
  MUX4ND0BWP U6814 ( .I0(\srf/regTable[4][0] ), .I1(\srf/regTable[5][0] ), 
        .I2(\srf/regTable[6][0] ), .I3(\srf/regTable[7][0] ), .S0(n4795), .S1(
        n4865), .ZN(n4565) );
  MUX2ND0BWP U6815 ( .I0(n4566), .I1(n4567), .S(n4915), .ZN(scalarData1[15])
         );
  MUX4ND0BWP U6816 ( .I0(\srf/regTable[0][15] ), .I1(\srf/regTable[1][15] ), 
        .I2(\srf/regTable[2][15] ), .I3(\srf/regTable[3][15] ), .S0(n4798), 
        .S1(n4868), .ZN(n4566) );
  MUX4ND0BWP U6817 ( .I0(\srf/regTable[4][15] ), .I1(\srf/regTable[5][15] ), 
        .I2(\srf/regTable[6][15] ), .I3(\srf/regTable[7][15] ), .S0(n4798), 
        .S1(n4868), .ZN(n4567) );
  MUX2ND0BWP U6818 ( .I0(n4568), .I1(n4569), .S(n4915), .ZN(scalarData1[14])
         );
  MUX4ND0BWP U6819 ( .I0(\srf/regTable[0][14] ), .I1(\srf/regTable[1][14] ), 
        .I2(\srf/regTable[2][14] ), .I3(\srf/regTable[3][14] ), .S0(n4798), 
        .S1(n4868), .ZN(n4568) );
  MUX4ND0BWP U6820 ( .I0(\srf/regTable[4][14] ), .I1(\srf/regTable[5][14] ), 
        .I2(\srf/regTable[6][14] ), .I3(\srf/regTable[7][14] ), .S0(n4798), 
        .S1(n4868), .ZN(n4569) );
  MUX2ND0BWP U6821 ( .I0(n4570), .I1(n4571), .S(n4915), .ZN(scalarData1[13])
         );
  MUX4ND0BWP U6822 ( .I0(\srf/regTable[0][13] ), .I1(\srf/regTable[1][13] ), 
        .I2(\srf/regTable[2][13] ), .I3(\srf/regTable[3][13] ), .S0(n4797), 
        .S1(n4867), .ZN(n4570) );
  MUX4ND0BWP U6823 ( .I0(\srf/regTable[4][13] ), .I1(\srf/regTable[5][13] ), 
        .I2(\srf/regTable[6][13] ), .I3(\srf/regTable[7][13] ), .S0(n4797), 
        .S1(n4867), .ZN(n4571) );
  MUX2ND0BWP U6824 ( .I0(n4572), .I1(n4573), .S(n4915), .ZN(scalarData1[12])
         );
  MUX4ND0BWP U6825 ( .I0(\srf/regTable[0][12] ), .I1(\srf/regTable[1][12] ), 
        .I2(\srf/regTable[2][12] ), .I3(\srf/regTable[3][12] ), .S0(n4797), 
        .S1(n4867), .ZN(n4572) );
  MUX4ND0BWP U6826 ( .I0(\srf/regTable[4][12] ), .I1(\srf/regTable[5][12] ), 
        .I2(\srf/regTable[6][12] ), .I3(\srf/regTable[7][12] ), .S0(n4797), 
        .S1(n4867), .ZN(n4573) );
  MUX2ND0BWP U6827 ( .I0(n4574), .I1(n4575), .S(n4915), .ZN(scalarData1[11])
         );
  MUX4ND0BWP U6828 ( .I0(\srf/regTable[0][11] ), .I1(\srf/regTable[1][11] ), 
        .I2(\srf/regTable[2][11] ), .I3(\srf/regTable[3][11] ), .S0(n4797), 
        .S1(n4867), .ZN(n4574) );
  MUX4ND0BWP U6829 ( .I0(\srf/regTable[4][11] ), .I1(\srf/regTable[5][11] ), 
        .I2(\srf/regTable[6][11] ), .I3(\srf/regTable[7][11] ), .S0(n4797), 
        .S1(n4867), .ZN(n4575) );
  MUX2ND0BWP U6830 ( .I0(n4576), .I1(n4577), .S(n4915), .ZN(scalarData1[10])
         );
  MUX4ND0BWP U6831 ( .I0(\srf/regTable[0][10] ), .I1(\srf/regTable[1][10] ), 
        .I2(\srf/regTable[2][10] ), .I3(\srf/regTable[3][10] ), .S0(n4797), 
        .S1(n4867), .ZN(n4576) );
  MUX4ND0BWP U6832 ( .I0(\srf/regTable[4][10] ), .I1(\srf/regTable[5][10] ), 
        .I2(\srf/regTable[6][10] ), .I3(\srf/regTable[7][10] ), .S0(n4797), 
        .S1(n4867), .ZN(n4577) );
  MUX2ND0BWP U6833 ( .I0(n4578), .I1(n4579), .S(n4915), .ZN(scalarData1[9]) );
  MUX4ND0BWP U6834 ( .I0(\srf/regTable[0][9] ), .I1(\srf/regTable[1][9] ), 
        .I2(\srf/regTable[2][9] ), .I3(\srf/regTable[3][9] ), .S0(n4797), .S1(
        n4867), .ZN(n4578) );
  MUX4ND0BWP U6835 ( .I0(\srf/regTable[4][9] ), .I1(\srf/regTable[5][9] ), 
        .I2(\srf/regTable[6][9] ), .I3(\srf/regTable[7][9] ), .S0(n4797), .S1(
        n4867), .ZN(n4579) );
  MUX2ND0BWP U6836 ( .I0(n4580), .I1(n4581), .S(n4915), .ZN(scalarData1[8]) );
  MUX4ND0BWP U6837 ( .I0(\srf/regTable[0][8] ), .I1(\srf/regTable[1][8] ), 
        .I2(\srf/regTable[2][8] ), .I3(\srf/regTable[3][8] ), .S0(n4797), .S1(
        n4867), .ZN(n4580) );
  MUX4ND0BWP U6838 ( .I0(\srf/regTable[4][8] ), .I1(\srf/regTable[5][8] ), 
        .I2(\srf/regTable[6][8] ), .I3(\srf/regTable[7][8] ), .S0(n4797), .S1(
        n4867), .ZN(n4581) );
  MUX2ND0BWP U6839 ( .I0(n4582), .I1(n4583), .S(n4914), .ZN(scalarData1[1]) );
  MUX4ND0BWP U6840 ( .I0(\srf/regTable[0][1] ), .I1(\srf/regTable[1][1] ), 
        .I2(\srf/regTable[2][1] ), .I3(\srf/regTable[3][1] ), .S0(n4795), .S1(
        n4865), .ZN(n4582) );
  MUX4ND0BWP U6841 ( .I0(\srf/regTable[4][1] ), .I1(\srf/regTable[5][1] ), 
        .I2(\srf/regTable[6][1] ), .I3(\srf/regTable[7][1] ), .S0(n4795), .S1(
        n4865), .ZN(n4583) );
  MUX2ND0BWP U6842 ( .I0(n4584), .I1(n4585), .S(n4914), .ZN(scalarData1[7]) );
  MUX4ND0BWP U6843 ( .I0(\srf/regTable[0][7] ), .I1(\srf/regTable[1][7] ), 
        .I2(\srf/regTable[2][7] ), .I3(\srf/regTable[3][7] ), .S0(n4796), .S1(
        n4866), .ZN(n4584) );
  MUX4ND0BWP U6844 ( .I0(\srf/regTable[4][7] ), .I1(\srf/regTable[5][7] ), 
        .I2(\srf/regTable[6][7] ), .I3(\srf/regTable[7][7] ), .S0(n4796), .S1(
        n4866), .ZN(n4585) );
  MUX2ND0BWP U6845 ( .I0(n4586), .I1(n4587), .S(n4914), .ZN(scalarData1[6]) );
  MUX4ND0BWP U6846 ( .I0(\srf/regTable[0][6] ), .I1(\srf/regTable[1][6] ), 
        .I2(\srf/regTable[2][6] ), .I3(\srf/regTable[3][6] ), .S0(n4796), .S1(
        n4866), .ZN(n4586) );
  MUX4ND0BWP U6847 ( .I0(\srf/regTable[4][6] ), .I1(\srf/regTable[5][6] ), 
        .I2(\srf/regTable[6][6] ), .I3(\srf/regTable[7][6] ), .S0(n4796), .S1(
        n4866), .ZN(n4587) );
  MUX2ND0BWP U6848 ( .I0(n4588), .I1(n4589), .S(n4914), .ZN(scalarData1[5]) );
  MUX4ND0BWP U6849 ( .I0(\srf/regTable[0][5] ), .I1(\srf/regTable[1][5] ), 
        .I2(\srf/regTable[2][5] ), .I3(\srf/regTable[3][5] ), .S0(n4796), .S1(
        n4866), .ZN(n4588) );
  MUX4ND0BWP U6850 ( .I0(\srf/regTable[4][5] ), .I1(\srf/regTable[5][5] ), 
        .I2(\srf/regTable[6][5] ), .I3(\srf/regTable[7][5] ), .S0(n4796), .S1(
        n4866), .ZN(n4589) );
  MUX2ND0BWP U6851 ( .I0(n4590), .I1(n4591), .S(n4914), .ZN(scalarData1[2]) );
  MUX4ND0BWP U6852 ( .I0(\srf/regTable[0][2] ), .I1(\srf/regTable[1][2] ), 
        .I2(\srf/regTable[2][2] ), .I3(\srf/regTable[3][2] ), .S0(n4796), .S1(
        n4866), .ZN(n4590) );
  MUX4ND0BWP U6853 ( .I0(\srf/regTable[4][2] ), .I1(\srf/regTable[5][2] ), 
        .I2(\srf/regTable[6][2] ), .I3(\srf/regTable[7][2] ), .S0(n4796), .S1(
        n4866), .ZN(n4591) );
  MUX2ND0BWP U6854 ( .I0(n4592), .I1(n4593), .S(n4914), .ZN(scalarData1[3]) );
  MUX4ND0BWP U6855 ( .I0(\srf/regTable[0][3] ), .I1(\srf/regTable[1][3] ), 
        .I2(\srf/regTable[2][3] ), .I3(\srf/regTable[3][3] ), .S0(n4796), .S1(
        n4866), .ZN(n4592) );
  MUX4ND0BWP U6856 ( .I0(\srf/regTable[4][3] ), .I1(\srf/regTable[5][3] ), 
        .I2(\srf/regTable[6][3] ), .I3(\srf/regTable[7][3] ), .S0(n4796), .S1(
        n4866), .ZN(n4593) );
  MUX2ND0BWP U6857 ( .I0(n4594), .I1(n4595), .S(n4914), .ZN(scalarData1[4]) );
  MUX4ND0BWP U6858 ( .I0(\srf/regTable[0][4] ), .I1(\srf/regTable[1][4] ), 
        .I2(\srf/regTable[2][4] ), .I3(\srf/regTable[3][4] ), .S0(n4796), .S1(
        n4866), .ZN(n4594) );
  MUX4ND0BWP U6859 ( .I0(\srf/regTable[4][4] ), .I1(\srf/regTable[5][4] ), 
        .I2(\srf/regTable[6][4] ), .I3(\srf/regTable[7][4] ), .S0(n4796), .S1(
        n4866), .ZN(n4595) );
  MUX2ND0BWP U6860 ( .I0(n4596), .I1(n4597), .S(n4893), .ZN(vectorData1[0]) );
  MUX4ND0BWP U6861 ( .I0(\vrf/regTable[0][0] ), .I1(\vrf/regTable[1][0] ), 
        .I2(\vrf/regTable[2][0] ), .I3(\vrf/regTable[3][0] ), .S0(n4753), .S1(
        n4823), .ZN(n4596) );
  MUX4ND0BWP U6862 ( .I0(\vrf/regTable[4][0] ), .I1(\vrf/regTable[5][0] ), 
        .I2(\vrf/regTable[6][0] ), .I3(\vrf/regTable[7][0] ), .S0(n4753), .S1(
        n4823), .ZN(n4597) );
  MUX2ND0BWP U6863 ( .I0(n4598), .I1(n4599), .S(n4894), .ZN(vectorData1[15])
         );
  MUX4ND0BWP U6864 ( .I0(\vrf/regTable[0][15] ), .I1(\vrf/regTable[1][15] ), 
        .I2(\vrf/regTable[2][15] ), .I3(\vrf/regTable[3][15] ), .S0(n4755), 
        .S1(n4825), .ZN(n4598) );
  MUX4ND0BWP U6865 ( .I0(\vrf/regTable[4][15] ), .I1(\vrf/regTable[5][15] ), 
        .I2(\vrf/regTable[6][15] ), .I3(\vrf/regTable[7][15] ), .S0(n4755), 
        .S1(n4825), .ZN(n4599) );
  MUX2ND0BWP U6866 ( .I0(n4600), .I1(n4601), .S(n4894), .ZN(vectorData1[14])
         );
  MUX4ND0BWP U6867 ( .I0(\vrf/regTable[0][14] ), .I1(\vrf/regTable[1][14] ), 
        .I2(\vrf/regTable[2][14] ), .I3(\vrf/regTable[3][14] ), .S0(n4755), 
        .S1(n4825), .ZN(n4600) );
  MUX4ND0BWP U6868 ( .I0(\vrf/regTable[4][14] ), .I1(\vrf/regTable[5][14] ), 
        .I2(\vrf/regTable[6][14] ), .I3(\vrf/regTable[7][14] ), .S0(n4755), 
        .S1(n4825), .ZN(n4601) );
  MUX2ND0BWP U6869 ( .I0(n4602), .I1(n4603), .S(n4894), .ZN(vectorData1[13])
         );
  MUX4ND0BWP U6870 ( .I0(\vrf/regTable[0][13] ), .I1(\vrf/regTable[1][13] ), 
        .I2(\vrf/regTable[2][13] ), .I3(\vrf/regTable[3][13] ), .S0(n4755), 
        .S1(n4825), .ZN(n4602) );
  MUX4ND0BWP U6871 ( .I0(\vrf/regTable[4][13] ), .I1(\vrf/regTable[5][13] ), 
        .I2(\vrf/regTable[6][13] ), .I3(\vrf/regTable[7][13] ), .S0(n4755), 
        .S1(n4825), .ZN(n4603) );
  MUX2ND0BWP U6872 ( .I0(n4604), .I1(n4605), .S(n4894), .ZN(vectorData1[12])
         );
  MUX4ND0BWP U6873 ( .I0(\vrf/regTable[0][12] ), .I1(\vrf/regTable[1][12] ), 
        .I2(\vrf/regTable[2][12] ), .I3(\vrf/regTable[3][12] ), .S0(n4755), 
        .S1(n4825), .ZN(n4604) );
  MUX4ND0BWP U6874 ( .I0(\vrf/regTable[4][12] ), .I1(\vrf/regTable[5][12] ), 
        .I2(\vrf/regTable[6][12] ), .I3(\vrf/regTable[7][12] ), .S0(n4755), 
        .S1(n4825), .ZN(n4605) );
  MUX2ND0BWP U6875 ( .I0(n4606), .I1(n4607), .S(n4893), .ZN(vectorData1[11])
         );
  MUX4ND0BWP U6876 ( .I0(\vrf/regTable[0][11] ), .I1(\vrf/regTable[1][11] ), 
        .I2(\vrf/regTable[2][11] ), .I3(\vrf/regTable[3][11] ), .S0(n4754), 
        .S1(n4824), .ZN(n4606) );
  MUX4ND0BWP U6877 ( .I0(\vrf/regTable[4][11] ), .I1(\vrf/regTable[5][11] ), 
        .I2(\vrf/regTable[6][11] ), .I3(\vrf/regTable[7][11] ), .S0(n4754), 
        .S1(n4824), .ZN(n4607) );
  MUX2ND0BWP U6878 ( .I0(n4608), .I1(n4609), .S(n4893), .ZN(vectorData1[10])
         );
  MUX4ND0BWP U6879 ( .I0(\vrf/regTable[0][10] ), .I1(\vrf/regTable[1][10] ), 
        .I2(\vrf/regTable[2][10] ), .I3(\vrf/regTable[3][10] ), .S0(n4754), 
        .S1(n4824), .ZN(n4608) );
  MUX4ND0BWP U6880 ( .I0(\vrf/regTable[4][10] ), .I1(\vrf/regTable[5][10] ), 
        .I2(\vrf/regTable[6][10] ), .I3(\vrf/regTable[7][10] ), .S0(n4754), 
        .S1(n4824), .ZN(n4609) );
  MUX2ND0BWP U6881 ( .I0(n4610), .I1(n4611), .S(n4893), .ZN(vectorData1[9]) );
  MUX4ND0BWP U6882 ( .I0(\vrf/regTable[0][9] ), .I1(\vrf/regTable[1][9] ), 
        .I2(\vrf/regTable[2][9] ), .I3(\vrf/regTable[3][9] ), .S0(n4754), .S1(
        n4824), .ZN(n4610) );
  MUX4ND0BWP U6883 ( .I0(\vrf/regTable[4][9] ), .I1(\vrf/regTable[5][9] ), 
        .I2(\vrf/regTable[6][9] ), .I3(\vrf/regTable[7][9] ), .S0(n4754), .S1(
        n4824), .ZN(n4611) );
  MUX2ND0BWP U6884 ( .I0(n4612), .I1(n4613), .S(n4893), .ZN(vectorData1[8]) );
  MUX4ND0BWP U6885 ( .I0(\vrf/regTable[0][8] ), .I1(\vrf/regTable[1][8] ), 
        .I2(\vrf/regTable[2][8] ), .I3(\vrf/regTable[3][8] ), .S0(n4754), .S1(
        n4824), .ZN(n4612) );
  MUX4ND0BWP U6886 ( .I0(\vrf/regTable[4][8] ), .I1(\vrf/regTable[5][8] ), 
        .I2(\vrf/regTable[6][8] ), .I3(\vrf/regTable[7][8] ), .S0(n4754), .S1(
        n4824), .ZN(n4613) );
  MUX2ND0BWP U6887 ( .I0(n4614), .I1(n4615), .S(n4893), .ZN(vectorData1[1]) );
  MUX4ND0BWP U6888 ( .I0(\vrf/regTable[0][1] ), .I1(\vrf/regTable[1][1] ), 
        .I2(\vrf/regTable[2][1] ), .I3(\vrf/regTable[3][1] ), .S0(n4753), .S1(
        n4823), .ZN(n4614) );
  MUX4ND0BWP U6889 ( .I0(\vrf/regTable[4][1] ), .I1(\vrf/regTable[5][1] ), 
        .I2(\vrf/regTable[6][1] ), .I3(\vrf/regTable[7][1] ), .S0(n4753), .S1(
        n4823), .ZN(n4615) );
  MUX2ND0BWP U6890 ( .I0(n4616), .I1(n4617), .S(n4893), .ZN(vectorData1[7]) );
  MUX4ND0BWP U6891 ( .I0(\vrf/regTable[0][7] ), .I1(\vrf/regTable[1][7] ), 
        .I2(\vrf/regTable[2][7] ), .I3(\vrf/regTable[3][7] ), .S0(n4754), .S1(
        n4824), .ZN(n4616) );
  MUX4ND0BWP U6892 ( .I0(\vrf/regTable[4][7] ), .I1(\vrf/regTable[5][7] ), 
        .I2(\vrf/regTable[6][7] ), .I3(\vrf/regTable[7][7] ), .S0(n4754), .S1(
        n4824), .ZN(n4617) );
  MUX2ND0BWP U6893 ( .I0(n4618), .I1(n4619), .S(n4893), .ZN(vectorData1[6]) );
  MUX4ND0BWP U6894 ( .I0(\vrf/regTable[0][6] ), .I1(\vrf/regTable[1][6] ), 
        .I2(\vrf/regTable[2][6] ), .I3(\vrf/regTable[3][6] ), .S0(n4754), .S1(
        n4824), .ZN(n4618) );
  MUX4ND0BWP U6895 ( .I0(\vrf/regTable[4][6] ), .I1(\vrf/regTable[5][6] ), 
        .I2(\vrf/regTable[6][6] ), .I3(\vrf/regTable[7][6] ), .S0(n4754), .S1(
        n4824), .ZN(n4619) );
  MUX2ND0BWP U6896 ( .I0(n4620), .I1(n4621), .S(n4893), .ZN(vectorData1[5]) );
  MUX4ND0BWP U6897 ( .I0(\vrf/regTable[0][5] ), .I1(\vrf/regTable[1][5] ), 
        .I2(\vrf/regTable[2][5] ), .I3(\vrf/regTable[3][5] ), .S0(n4753), .S1(
        n4823), .ZN(n4620) );
  MUX4ND0BWP U6898 ( .I0(\vrf/regTable[4][5] ), .I1(\vrf/regTable[5][5] ), 
        .I2(\vrf/regTable[6][5] ), .I3(\vrf/regTable[7][5] ), .S0(n4753), .S1(
        n4823), .ZN(n4621) );
  MUX2ND0BWP U6899 ( .I0(n4622), .I1(n4623), .S(n4893), .ZN(vectorData1[2]) );
  MUX4ND0BWP U6900 ( .I0(\vrf/regTable[0][2] ), .I1(\vrf/regTable[1][2] ), 
        .I2(\vrf/regTable[2][2] ), .I3(\vrf/regTable[3][2] ), .S0(n4753), .S1(
        n4823), .ZN(n4622) );
  MUX4ND0BWP U6901 ( .I0(\vrf/regTable[4][2] ), .I1(\vrf/regTable[5][2] ), 
        .I2(\vrf/regTable[6][2] ), .I3(\vrf/regTable[7][2] ), .S0(n4753), .S1(
        n4823), .ZN(n4623) );
  MUX2ND0BWP U6902 ( .I0(n4624), .I1(n4625), .S(n4893), .ZN(vectorData1[3]) );
  MUX4ND0BWP U6903 ( .I0(\vrf/regTable[0][3] ), .I1(\vrf/regTable[1][3] ), 
        .I2(\vrf/regTable[2][3] ), .I3(\vrf/regTable[3][3] ), .S0(n4753), .S1(
        n4823), .ZN(n4624) );
  MUX4ND0BWP U6904 ( .I0(\vrf/regTable[4][3] ), .I1(\vrf/regTable[5][3] ), 
        .I2(\vrf/regTable[6][3] ), .I3(\vrf/regTable[7][3] ), .S0(n4753), .S1(
        n4823), .ZN(n4625) );
  MUX2ND0BWP U6905 ( .I0(n4626), .I1(n4627), .S(n4893), .ZN(vectorData1[4]) );
  MUX4ND0BWP U6906 ( .I0(\vrf/regTable[0][4] ), .I1(\vrf/regTable[1][4] ), 
        .I2(\vrf/regTable[2][4] ), .I3(\vrf/regTable[3][4] ), .S0(n4753), .S1(
        n4823), .ZN(n4626) );
  MUX4ND0BWP U6907 ( .I0(\vrf/regTable[4][4] ), .I1(\vrf/regTable[5][4] ), 
        .I2(\vrf/regTable[6][4] ), .I3(\vrf/regTable[7][4] ), .S0(n4753), .S1(
        n4823), .ZN(n4627) );
  CKBD1BWP U6908 ( .I(\vrf/N11 ), .Z(n4927) );
  OR2XD1BWP U6909 ( .A1(func[3]), .A2(n4628), .Z(n5468) );
  MUX2ND0BWP U6910 ( .I0(op1[15]), .I1(op2[7]), .S(func[0]), .ZN(n4628) );
  TIELBWP U6911 ( .ZN(\*Logic0* ) );
  TIEHBWP U6912 ( .Z(\alu/*Logic1* ) );
  INR2D0BWP U6913 ( .A1(n7371), .B1(n4639), .ZN(\vrf/N99 ) );
  INR2D0BWP U6914 ( .A1(n7372), .B1(n4639), .ZN(\vrf/N98 ) );
  INR2D0BWP U6915 ( .A1(n7373), .B1(n4638), .ZN(\vrf/N97 ) );
  INR2D0BWP U6916 ( .A1(n7374), .B1(n4638), .ZN(\vrf/N96 ) );
  INR2D0BWP U6917 ( .A1(n7375), .B1(n4638), .ZN(\vrf/N95 ) );
  INR2D0BWP U6918 ( .A1(n7376), .B1(n4638), .ZN(\vrf/N94 ) );
  INR2D0BWP U6919 ( .A1(n7377), .B1(n4638), .ZN(\vrf/N93 ) );
  INR2D0BWP U6920 ( .A1(n7378), .B1(n4638), .ZN(\vrf/N92 ) );
  INR2D0BWP U6921 ( .A1(n7379), .B1(n4638), .ZN(\vrf/N91 ) );
  INR2D0BWP U6922 ( .A1(n7380), .B1(n4638), .ZN(\vrf/N90 ) );
  OAI22D0BWP U6923 ( .A1(n5525), .A2(n5526), .B1(n5527), .B2(n5528), .ZN(
        \vrf/N9 ) );
  CKND0BWP U6924 ( .I(instrIn[6]), .ZN(n5528) );
  INR2D0BWP U6925 ( .A1(n7381), .B1(n4638), .ZN(\vrf/N89 ) );
  INR2D0BWP U6926 ( .A1(n7382), .B1(n4638), .ZN(\vrf/N88 ) );
  INR2D0BWP U6927 ( .A1(n7383), .B1(n4638), .ZN(\vrf/N87 ) );
  INR2D0BWP U6928 ( .A1(n7384), .B1(n4638), .ZN(\vrf/N86 ) );
  INR2D0BWP U6929 ( .A1(n7385), .B1(n4638), .ZN(\vrf/N85 ) );
  INR2D0BWP U6930 ( .A1(n7386), .B1(n4637), .ZN(\vrf/N84 ) );
  INR2D0BWP U6931 ( .A1(n7387), .B1(n4637), .ZN(\vrf/N83 ) );
  INR2D0BWP U6932 ( .A1(n7388), .B1(n4637), .ZN(\vrf/N82 ) );
  INR2D0BWP U6933 ( .A1(n7389), .B1(n4637), .ZN(\vrf/N81 ) );
  INR2D0BWP U6934 ( .A1(n7390), .B1(n4637), .ZN(\vrf/N80 ) );
  INR2D0BWP U6935 ( .A1(n7391), .B1(n4637), .ZN(\vrf/N79 ) );
  INR2D0BWP U6936 ( .A1(n7392), .B1(n4637), .ZN(\vrf/N78 ) );
  INR2D0BWP U6937 ( .A1(n7393), .B1(n4637), .ZN(\vrf/N77 ) );
  INR2D0BWP U6938 ( .A1(n7394), .B1(n4637), .ZN(\vrf/N76 ) );
  INR2D0BWP U6939 ( .A1(n7395), .B1(n4637), .ZN(\vrf/N75 ) );
  INR2D0BWP U6940 ( .A1(n7396), .B1(n4637), .ZN(\vrf/N74 ) );
  INR2D0BWP U6941 ( .A1(n7397), .B1(n4637), .ZN(\vrf/N73 ) );
  INR2D0BWP U6942 ( .A1(n7398), .B1(n4637), .ZN(\vrf/N72 ) );
  INR2D0BWP U6943 ( .A1(n7399), .B1(n4636), .ZN(\vrf/N71 ) );
  INR2D0BWP U6944 ( .A1(n7400), .B1(n4636), .ZN(\vrf/N70 ) );
  INR2D0BWP U6945 ( .A1(n7401), .B1(n4636), .ZN(\vrf/N69 ) );
  INR2D0BWP U6946 ( .A1(n7402), .B1(n4636), .ZN(\vrf/N68 ) );
  INR2D0BWP U6947 ( .A1(n7403), .B1(n4636), .ZN(\vrf/N67 ) );
  INR2D0BWP U6948 ( .A1(n7404), .B1(n4636), .ZN(\vrf/N66 ) );
  INR2D0BWP U6949 ( .A1(n7405), .B1(n4636), .ZN(\vrf/N65 ) );
  INR2D0BWP U6950 ( .A1(n7406), .B1(n4636), .ZN(\vrf/N64 ) );
  INR2D0BWP U6951 ( .A1(n7407), .B1(n4636), .ZN(\vrf/N63 ) );
  INR2D0BWP U6952 ( .A1(n7408), .B1(n4636), .ZN(\vrf/N62 ) );
  INR2D0BWP U6953 ( .A1(n7409), .B1(n4636), .ZN(\vrf/N61 ) );
  INR2D0BWP U6954 ( .A1(n7410), .B1(n4636), .ZN(\vrf/N60 ) );
  INR2D0BWP U6955 ( .A1(n7411), .B1(n4636), .ZN(\vrf/N59 ) );
  INR2D0BWP U6956 ( .A1(n7412), .B1(n4635), .ZN(\vrf/N58 ) );
  INR2D0BWP U6957 ( .A1(n7413), .B1(n4635), .ZN(\vrf/N57 ) );
  INR2D0BWP U6958 ( .A1(n7414), .B1(n4635), .ZN(\vrf/N56 ) );
  INR2D0BWP U6959 ( .A1(n7415), .B1(n4635), .ZN(\vrf/N55 ) );
  INR2D0BWP U6960 ( .A1(n7416), .B1(n4635), .ZN(\vrf/N54 ) );
  INR2D0BWP U6961 ( .A1(n7417), .B1(n4635), .ZN(\vrf/N53 ) );
  INR2D0BWP U6962 ( .A1(n7418), .B1(n4635), .ZN(\vrf/N52 ) );
  INR2D0BWP U6963 ( .A1(n7419), .B1(n4635), .ZN(\vrf/N51 ) );
  INR2D0BWP U6964 ( .A1(n7420), .B1(n4635), .ZN(\vrf/N50 ) );
  INR2D0BWP U6965 ( .A1(n7421), .B1(n4635), .ZN(\vrf/N49 ) );
  INR2D0BWP U6966 ( .A1(n7422), .B1(n4635), .ZN(\vrf/N48 ) );
  INR2D0BWP U6967 ( .A1(n7423), .B1(n4635), .ZN(\vrf/N47 ) );
  INR2D0BWP U6968 ( .A1(n7424), .B1(n4635), .ZN(\vrf/N46 ) );
  INR2D0BWP U6969 ( .A1(n7425), .B1(n4634), .ZN(\vrf/N45 ) );
  INR2D0BWP U6970 ( .A1(n7426), .B1(n4634), .ZN(\vrf/N44 ) );
  INR2D0BWP U6971 ( .A1(n7427), .B1(n4634), .ZN(\vrf/N43 ) );
  INR2D0BWP U6972 ( .A1(n7428), .B1(n4634), .ZN(\vrf/N42 ) );
  INR2D0BWP U6973 ( .A1(n7429), .B1(n4634), .ZN(\vrf/N41 ) );
  INR2D0BWP U6974 ( .A1(n7430), .B1(n4634), .ZN(\vrf/N40 ) );
  INR2D0BWP U6975 ( .A1(n7431), .B1(n4634), .ZN(\vrf/N39 ) );
  INR2D0BWP U6976 ( .A1(n7432), .B1(n4634), .ZN(\vrf/N38 ) );
  INR2D0BWP U6977 ( .A1(n7433), .B1(n4634), .ZN(\vrf/N37 ) );
  INR2D0BWP U6978 ( .A1(n7434), .B1(n4634), .ZN(\vrf/N36 ) );
  INR2D0BWP U6979 ( .A1(n7435), .B1(n4634), .ZN(\vrf/N35 ) );
  NR2D0BWP U6980 ( .A1(n4629), .A2(n3419), .ZN(\vrf/N34 ) );
  NR2D0BWP U6981 ( .A1(n4630), .A2(n3403), .ZN(\vrf/N33 ) );
  NR2D0BWP U6982 ( .A1(n4630), .A2(n3404), .ZN(\vrf/N32 ) );
  NR2D0BWP U6983 ( .A1(n4630), .A2(n3405), .ZN(\vrf/N31 ) );
  NR2D0BWP U6984 ( .A1(n4630), .A2(n3406), .ZN(\vrf/N30 ) );
  OAI21D0BWP U6985 ( .A1(n5529), .A2(n5530), .B(n7436), .ZN(\vrf/N296 ) );
  OAI21D0BWP U6986 ( .A1(n5530), .A2(n5531), .B(n7436), .ZN(\vrf/N293 ) );
  OAI21D0BWP U6987 ( .A1(n5529), .A2(n5532), .B(n7436), .ZN(\vrf/N290 ) );
  NR2D0BWP U6988 ( .A1(n4629), .A2(n3407), .ZN(\vrf/N29 ) );
  OAI21D0BWP U6989 ( .A1(n5531), .A2(n5532), .B(n7436), .ZN(\vrf/N287 ) );
  OAI21D0BWP U6990 ( .A1(n5529), .A2(n5533), .B(n7436), .ZN(\vrf/N284 ) );
  OAI21D0BWP U6991 ( .A1(n5531), .A2(n5533), .B(n7436), .ZN(\vrf/N281 ) );
  NR2D0BWP U6992 ( .A1(n4629), .A2(n3408), .ZN(\vrf/N28 ) );
  OAI21D0BWP U6993 ( .A1(n5529), .A2(n5534), .B(n7436), .ZN(\vrf/N278 ) );
  CKND2D0BWP U6994 ( .A1(n5535), .A2(n7437), .ZN(n5529) );
  INR2D0BWP U6995 ( .A1(n7197), .B1(n4633), .ZN(\vrf/N275 ) );
  INR2D0BWP U6996 ( .A1(n7198), .B1(n4633), .ZN(\vrf/N274 ) );
  INR2D0BWP U6997 ( .A1(n7199), .B1(n4633), .ZN(\vrf/N273 ) );
  INR2D0BWP U6998 ( .A1(n7200), .B1(n4633), .ZN(\vrf/N272 ) );
  INR2D0BWP U6999 ( .A1(n7201), .B1(n4633), .ZN(\vrf/N271 ) );
  INR2D0BWP U7000 ( .A1(n7202), .B1(n4633), .ZN(\vrf/N270 ) );
  NR2D0BWP U7001 ( .A1(n4630), .A2(n3409), .ZN(\vrf/N27 ) );
  INR2D0BWP U7002 ( .A1(n7203), .B1(n4633), .ZN(\vrf/N269 ) );
  INR2D0BWP U7003 ( .A1(n7204), .B1(n4633), .ZN(\vrf/N268 ) );
  INR2D0BWP U7004 ( .A1(n7205), .B1(n4632), .ZN(\vrf/N267 ) );
  INR2D0BWP U7005 ( .A1(n7206), .B1(n4633), .ZN(\vrf/N266 ) );
  INR2D0BWP U7006 ( .A1(n7207), .B1(n4632), .ZN(\vrf/N265 ) );
  INR2D0BWP U7007 ( .A1(n7208), .B1(n4633), .ZN(\vrf/N264 ) );
  INR2D0BWP U7008 ( .A1(n7209), .B1(n4632), .ZN(\vrf/N263 ) );
  INR2D0BWP U7009 ( .A1(n7210), .B1(n4633), .ZN(\vrf/N262 ) );
  INR2D0BWP U7010 ( .A1(n7211), .B1(n4632), .ZN(\vrf/N261 ) );
  INR2D0BWP U7011 ( .A1(n7212), .B1(n4632), .ZN(\vrf/N260 ) );
  NR2D0BWP U7012 ( .A1(n4629), .A2(n3410), .ZN(\vrf/N26 ) );
  INR2D0BWP U7013 ( .A1(n7213), .B1(n4632), .ZN(\vrf/N259 ) );
  INR2D0BWP U7014 ( .A1(n7214), .B1(n4632), .ZN(\vrf/N258 ) );
  INR2D0BWP U7015 ( .A1(n7215), .B1(n4634), .ZN(\vrf/N257 ) );
  INR2D0BWP U7016 ( .A1(n7216), .B1(n4633), .ZN(\vrf/N256 ) );
  INR2D0BWP U7017 ( .A1(n7217), .B1(n4631), .ZN(\vrf/N255 ) );
  INR2D0BWP U7018 ( .A1(n7218), .B1(n4632), .ZN(\vrf/N254 ) );
  INR2D0BWP U7019 ( .A1(n7219), .B1(n4631), .ZN(\vrf/N253 ) );
  INR2D0BWP U7020 ( .A1(n7220), .B1(n4632), .ZN(\vrf/N252 ) );
  INR2D0BWP U7021 ( .A1(n7221), .B1(n4632), .ZN(\vrf/N251 ) );
  INR2D0BWP U7022 ( .A1(n7222), .B1(n4631), .ZN(\vrf/N250 ) );
  NR2D0BWP U7023 ( .A1(n4629), .A2(n3411), .ZN(\vrf/N25 ) );
  INR2D0BWP U7024 ( .A1(n7223), .B1(n4633), .ZN(\vrf/N249 ) );
  INR2D0BWP U7025 ( .A1(n7224), .B1(n4632), .ZN(\vrf/N248 ) );
  INR2D0BWP U7026 ( .A1(n7225), .B1(n4631), .ZN(\vrf/N247 ) );
  INR2D0BWP U7027 ( .A1(n7226), .B1(n4631), .ZN(\vrf/N246 ) );
  INR2D0BWP U7028 ( .A1(n7227), .B1(n4630), .ZN(\vrf/N245 ) );
  INR2D0BWP U7029 ( .A1(n7228), .B1(n4631), .ZN(\vrf/N244 ) );
  INR2D0BWP U7030 ( .A1(n7229), .B1(n4631), .ZN(\vrf/N243 ) );
  INR2D0BWP U7031 ( .A1(n7230), .B1(n4631), .ZN(\vrf/N242 ) );
  INR2D0BWP U7032 ( .A1(n7231), .B1(n4631), .ZN(\vrf/N241 ) );
  INR2D0BWP U7033 ( .A1(n7232), .B1(n4630), .ZN(\vrf/N240 ) );
  NR2D0BWP U7034 ( .A1(n4629), .A2(n3412), .ZN(\vrf/N24 ) );
  INR2D0BWP U7035 ( .A1(n7233), .B1(n4630), .ZN(\vrf/N239 ) );
  INR2D0BWP U7036 ( .A1(n7234), .B1(n4632), .ZN(\vrf/N238 ) );
  INR2D0BWP U7037 ( .A1(n7235), .B1(n4630), .ZN(\vrf/N237 ) );
  INR2D0BWP U7038 ( .A1(n7236), .B1(n4631), .ZN(\vrf/N236 ) );
  INR2D0BWP U7039 ( .A1(n7237), .B1(n4632), .ZN(\vrf/N235 ) );
  INR2D0BWP U7040 ( .A1(n7238), .B1(n4631), .ZN(\vrf/N234 ) );
  INR2D0BWP U7041 ( .A1(n7239), .B1(n4631), .ZN(\vrf/N233 ) );
  INR2D0BWP U7042 ( .A1(n7240), .B1(n4630), .ZN(\vrf/N232 ) );
  INR2D0BWP U7043 ( .A1(n7241), .B1(n4630), .ZN(\vrf/N231 ) );
  INR2D0BWP U7044 ( .A1(n7242), .B1(n4630), .ZN(\vrf/N230 ) );
  NR2D0BWP U7045 ( .A1(n4629), .A2(n3413), .ZN(\vrf/N23 ) );
  INR2D0BWP U7046 ( .A1(n7243), .B1(n4630), .ZN(\vrf/N229 ) );
  INR2D0BWP U7047 ( .A1(n7244), .B1(n4634), .ZN(\vrf/N228 ) );
  INR2D0BWP U7048 ( .A1(n7245), .B1(n4648), .ZN(\vrf/N227 ) );
  INR2D0BWP U7049 ( .A1(n7246), .B1(n4648), .ZN(\vrf/N226 ) );
  INR2D0BWP U7050 ( .A1(n7247), .B1(n4648), .ZN(\vrf/N225 ) );
  INR2D0BWP U7051 ( .A1(n7248), .B1(n4648), .ZN(\vrf/N224 ) );
  INR2D0BWP U7052 ( .A1(n7249), .B1(n4648), .ZN(\vrf/N223 ) );
  INR2D0BWP U7053 ( .A1(n7250), .B1(n4648), .ZN(\vrf/N222 ) );
  INR2D0BWP U7054 ( .A1(n7251), .B1(n4648), .ZN(\vrf/N221 ) );
  INR2D0BWP U7055 ( .A1(n7252), .B1(n4648), .ZN(\vrf/N220 ) );
  NR2D0BWP U7056 ( .A1(n4629), .A2(n3414), .ZN(\vrf/N22 ) );
  INR2D0BWP U7057 ( .A1(n7253), .B1(n4648), .ZN(\vrf/N219 ) );
  INR2D0BWP U7058 ( .A1(n7254), .B1(n4648), .ZN(\vrf/N218 ) );
  OAI21D0BWP U7059 ( .A1(n5531), .A2(n5534), .B(n7436), .ZN(\vrf/N217 ) );
  CKND2D0BWP U7060 ( .A1(n5535), .A2(\srf/N15 ), .ZN(n5531) );
  INR2D0BWP U7061 ( .A1(n7255), .B1(n4647), .ZN(\vrf/N216 ) );
  INR2D0BWP U7062 ( .A1(n7256), .B1(n4647), .ZN(\vrf/N215 ) );
  INR2D0BWP U7063 ( .A1(n7257), .B1(n4647), .ZN(\vrf/N214 ) );
  INR2D0BWP U7064 ( .A1(n7258), .B1(n4647), .ZN(\vrf/N213 ) );
  INR2D0BWP U7065 ( .A1(n7259), .B1(n4647), .ZN(\vrf/N212 ) );
  INR2D0BWP U7066 ( .A1(n7260), .B1(n4647), .ZN(\vrf/N211 ) );
  INR2D0BWP U7067 ( .A1(n7261), .B1(n4647), .ZN(\vrf/N210 ) );
  NR2D0BWP U7068 ( .A1(n4629), .A2(n3415), .ZN(\vrf/N21 ) );
  INR2D0BWP U7069 ( .A1(n7262), .B1(n4647), .ZN(\vrf/N209 ) );
  INR2D0BWP U7070 ( .A1(n7263), .B1(n4647), .ZN(\vrf/N208 ) );
  INR2D0BWP U7071 ( .A1(n7264), .B1(n4647), .ZN(\vrf/N207 ) );
  INR2D0BWP U7072 ( .A1(n7265), .B1(n4647), .ZN(\vrf/N206 ) );
  INR2D0BWP U7073 ( .A1(n7266), .B1(n4647), .ZN(\vrf/N205 ) );
  INR2D0BWP U7074 ( .A1(n7267), .B1(n4647), .ZN(\vrf/N204 ) );
  INR2D0BWP U7075 ( .A1(n7268), .B1(n4646), .ZN(\vrf/N203 ) );
  INR2D0BWP U7076 ( .A1(n7269), .B1(n4646), .ZN(\vrf/N202 ) );
  INR2D0BWP U7077 ( .A1(n7270), .B1(n4646), .ZN(\vrf/N201 ) );
  INR2D0BWP U7078 ( .A1(n7271), .B1(n4646), .ZN(\vrf/N200 ) );
  NR2D0BWP U7079 ( .A1(n4629), .A2(n3416), .ZN(\vrf/N20 ) );
  INR2D0BWP U7080 ( .A1(n7272), .B1(n4646), .ZN(\vrf/N199 ) );
  INR2D0BWP U7081 ( .A1(n7273), .B1(n4646), .ZN(\vrf/N198 ) );
  INR2D0BWP U7082 ( .A1(n7274), .B1(n4646), .ZN(\vrf/N197 ) );
  INR2D0BWP U7083 ( .A1(n7275), .B1(n4646), .ZN(\vrf/N196 ) );
  INR2D0BWP U7084 ( .A1(n7276), .B1(n4646), .ZN(\vrf/N195 ) );
  INR2D0BWP U7085 ( .A1(n7277), .B1(n4646), .ZN(\vrf/N194 ) );
  INR2D0BWP U7086 ( .A1(n7278), .B1(n4646), .ZN(\vrf/N193 ) );
  INR2D0BWP U7087 ( .A1(n7279), .B1(n4646), .ZN(\vrf/N192 ) );
  INR2D0BWP U7088 ( .A1(n7280), .B1(n4646), .ZN(\vrf/N191 ) );
  INR2D0BWP U7089 ( .A1(n7281), .B1(n4645), .ZN(\vrf/N190 ) );
  NR2D0BWP U7090 ( .A1(n4629), .A2(n3417), .ZN(\vrf/N19 ) );
  INR2D0BWP U7091 ( .A1(n7282), .B1(n4645), .ZN(\vrf/N189 ) );
  INR2D0BWP U7092 ( .A1(n7283), .B1(n4645), .ZN(\vrf/N188 ) );
  INR2D0BWP U7093 ( .A1(n7284), .B1(n4645), .ZN(\vrf/N187 ) );
  INR2D0BWP U7094 ( .A1(n7285), .B1(n4645), .ZN(\vrf/N186 ) );
  INR2D0BWP U7095 ( .A1(n7286), .B1(n4645), .ZN(\vrf/N185 ) );
  INR2D0BWP U7096 ( .A1(n7287), .B1(n4645), .ZN(\vrf/N184 ) );
  INR2D0BWP U7097 ( .A1(n7288), .B1(n4645), .ZN(\vrf/N183 ) );
  INR2D0BWP U7098 ( .A1(n7289), .B1(n4645), .ZN(\vrf/N182 ) );
  INR2D0BWP U7099 ( .A1(n7290), .B1(n4645), .ZN(\vrf/N181 ) );
  INR2D0BWP U7100 ( .A1(n7291), .B1(n4645), .ZN(\vrf/N180 ) );
  NR2D0BWP U7101 ( .A1(n4629), .A2(n3418), .ZN(\vrf/N18 ) );
  INR2D0BWP U7102 ( .A1(n7292), .B1(n4645), .ZN(\vrf/N179 ) );
  INR2D0BWP U7103 ( .A1(n7293), .B1(n4645), .ZN(\vrf/N178 ) );
  INR2D0BWP U7104 ( .A1(n7294), .B1(n4644), .ZN(\vrf/N177 ) );
  INR2D0BWP U7105 ( .A1(n7295), .B1(n4644), .ZN(\vrf/N176 ) );
  INR2D0BWP U7106 ( .A1(n7296), .B1(n4644), .ZN(\vrf/N175 ) );
  INR2D0BWP U7107 ( .A1(n7297), .B1(n4644), .ZN(\vrf/N174 ) );
  INR2D0BWP U7108 ( .A1(n7298), .B1(n4644), .ZN(\vrf/N173 ) );
  INR2D0BWP U7109 ( .A1(n7299), .B1(n4644), .ZN(\vrf/N172 ) );
  INR2D0BWP U7110 ( .A1(n7300), .B1(n4644), .ZN(\vrf/N171 ) );
  INR2D0BWP U7111 ( .A1(n7301), .B1(n4644), .ZN(\vrf/N170 ) );
  INR2D0BWP U7112 ( .A1(n7302), .B1(n4644), .ZN(\vrf/N169 ) );
  INR2D0BWP U7113 ( .A1(n7303), .B1(n4644), .ZN(\vrf/N168 ) );
  INR2D0BWP U7114 ( .A1(n7304), .B1(n4644), .ZN(\vrf/N167 ) );
  INR2D0BWP U7115 ( .A1(n7305), .B1(n4644), .ZN(\vrf/N166 ) );
  INR2D0BWP U7116 ( .A1(n7306), .B1(n4644), .ZN(\vrf/N165 ) );
  INR2D0BWP U7117 ( .A1(n7307), .B1(n4643), .ZN(\vrf/N164 ) );
  INR2D0BWP U7118 ( .A1(n7308), .B1(n4643), .ZN(\vrf/N163 ) );
  INR2D0BWP U7119 ( .A1(n7309), .B1(n4643), .ZN(\vrf/N162 ) );
  INR2D0BWP U7120 ( .A1(n7310), .B1(n4643), .ZN(\vrf/N161 ) );
  INR2D0BWP U7121 ( .A1(n7311), .B1(n4643), .ZN(\vrf/N160 ) );
  INR2D0BWP U7122 ( .A1(n7312), .B1(n4643), .ZN(\vrf/N159 ) );
  INR2D0BWP U7123 ( .A1(n7313), .B1(n4643), .ZN(\vrf/N158 ) );
  INR2D0BWP U7124 ( .A1(n7314), .B1(n4643), .ZN(\vrf/N157 ) );
  INR2D0BWP U7125 ( .A1(n7315), .B1(n4643), .ZN(\vrf/N156 ) );
  INR2D0BWP U7126 ( .A1(n7316), .B1(n4643), .ZN(\vrf/N155 ) );
  INR2D0BWP U7127 ( .A1(n7317), .B1(n4643), .ZN(\vrf/N154 ) );
  INR2D0BWP U7128 ( .A1(n7318), .B1(n4643), .ZN(\vrf/N153 ) );
  INR2D0BWP U7129 ( .A1(n7319), .B1(n4642), .ZN(\vrf/N152 ) );
  INR2D0BWP U7130 ( .A1(n7320), .B1(n4642), .ZN(\vrf/N151 ) );
  INR2D0BWP U7131 ( .A1(n7321), .B1(n4642), .ZN(\vrf/N150 ) );
  INR2D0BWP U7132 ( .A1(n7322), .B1(n4642), .ZN(\vrf/N149 ) );
  INR2D0BWP U7133 ( .A1(n7323), .B1(n4642), .ZN(\vrf/N148 ) );
  INR2D0BWP U7134 ( .A1(n7324), .B1(n4642), .ZN(\vrf/N147 ) );
  INR2D0BWP U7135 ( .A1(n7325), .B1(n4642), .ZN(\vrf/N146 ) );
  INR2D0BWP U7136 ( .A1(n7326), .B1(n4642), .ZN(\vrf/N145 ) );
  INR2D0BWP U7137 ( .A1(n7327), .B1(n4642), .ZN(\vrf/N144 ) );
  INR2D0BWP U7138 ( .A1(n7328), .B1(n4642), .ZN(\vrf/N143 ) );
  INR2D0BWP U7139 ( .A1(n7329), .B1(n4642), .ZN(\vrf/N142 ) );
  INR2D0BWP U7140 ( .A1(n7330), .B1(n4642), .ZN(\vrf/N141 ) );
  INR2D0BWP U7141 ( .A1(n7331), .B1(n4642), .ZN(\vrf/N140 ) );
  OAI22D0BWP U7142 ( .A1(n5536), .A2(n5537), .B1(n5538), .B2(n5539), .ZN(
        \vrf/N14 ) );
  INR2D0BWP U7143 ( .A1(n7332), .B1(n4641), .ZN(\vrf/N139 ) );
  INR2D0BWP U7144 ( .A1(n7333), .B1(n4641), .ZN(\vrf/N138 ) );
  INR2D0BWP U7145 ( .A1(n7334), .B1(n4641), .ZN(\vrf/N137 ) );
  INR2D0BWP U7146 ( .A1(n7335), .B1(n4641), .ZN(\vrf/N136 ) );
  INR2D0BWP U7147 ( .A1(n7336), .B1(n4641), .ZN(\vrf/N135 ) );
  INR2D0BWP U7148 ( .A1(n7337), .B1(n4641), .ZN(\vrf/N134 ) );
  INR2D0BWP U7149 ( .A1(n7338), .B1(n4641), .ZN(\vrf/N133 ) );
  INR2D0BWP U7150 ( .A1(n7339), .B1(n4641), .ZN(\vrf/N132 ) );
  INR2D0BWP U7151 ( .A1(n7340), .B1(n4641), .ZN(\vrf/N131 ) );
  INR2D0BWP U7152 ( .A1(n7341), .B1(n4641), .ZN(\vrf/N130 ) );
  OAI22D0BWP U7153 ( .A1(n5536), .A2(n5540), .B1(n5538), .B2(n5541), .ZN(
        \vrf/N13 ) );
  INR2D0BWP U7154 ( .A1(n7342), .B1(n4641), .ZN(\vrf/N129 ) );
  INR2D0BWP U7155 ( .A1(n7343), .B1(n4641), .ZN(\vrf/N128 ) );
  INR2D0BWP U7156 ( .A1(n7344), .B1(n4641), .ZN(\vrf/N127 ) );
  INR2D0BWP U7157 ( .A1(n7345), .B1(n4640), .ZN(\vrf/N126 ) );
  INR2D0BWP U7158 ( .A1(n7346), .B1(n4640), .ZN(\vrf/N125 ) );
  INR2D0BWP U7159 ( .A1(n7347), .B1(n4640), .ZN(\vrf/N124 ) );
  INR2D0BWP U7160 ( .A1(n7348), .B1(n4640), .ZN(\vrf/N123 ) );
  INR2D0BWP U7161 ( .A1(n7349), .B1(n4640), .ZN(\vrf/N122 ) );
  INR2D0BWP U7162 ( .A1(n7350), .B1(n4640), .ZN(\vrf/N121 ) );
  INR2D0BWP U7163 ( .A1(n7351), .B1(n4640), .ZN(\vrf/N120 ) );
  OAI22D0BWP U7164 ( .A1(n5536), .A2(n5542), .B1(n5526), .B2(n5538), .ZN(
        \vrf/N12 ) );
  INR2D0BWP U7165 ( .A1(n7352), .B1(n4640), .ZN(\vrf/N119 ) );
  INR2D0BWP U7166 ( .A1(n7353), .B1(n4640), .ZN(\vrf/N118 ) );
  INR2D0BWP U7167 ( .A1(n7354), .B1(n4640), .ZN(\vrf/N116 ) );
  INR2D0BWP U7168 ( .A1(n7355), .B1(n4640), .ZN(\vrf/N115 ) );
  INR2D0BWP U7169 ( .A1(n7356), .B1(n4640), .ZN(\vrf/N114 ) );
  INR2D0BWP U7170 ( .A1(n7357), .B1(n4640), .ZN(\vrf/N113 ) );
  INR2D0BWP U7171 ( .A1(n7358), .B1(n4639), .ZN(\vrf/N112 ) );
  INR2D0BWP U7172 ( .A1(n7359), .B1(n4639), .ZN(\vrf/N111 ) );
  INR2D0BWP U7173 ( .A1(n7360), .B1(n4639), .ZN(\vrf/N110 ) );
  OAI22D0BWP U7174 ( .A1(n5525), .A2(n5539), .B1(n5527), .B2(n5543), .ZN(
        \vrf/N11 ) );
  CKND0BWP U7175 ( .I(instrIn[8]), .ZN(n5543) );
  INR2D0BWP U7176 ( .A1(n7361), .B1(n4639), .ZN(\vrf/N109 ) );
  INR2D0BWP U7177 ( .A1(n7362), .B1(n4639), .ZN(\vrf/N108 ) );
  INR2D0BWP U7178 ( .A1(n7363), .B1(n4639), .ZN(\vrf/N107 ) );
  INR2D0BWP U7179 ( .A1(n7364), .B1(n4639), .ZN(\vrf/N106 ) );
  INR2D0BWP U7180 ( .A1(n7365), .B1(n4639), .ZN(\vrf/N105 ) );
  INR2D0BWP U7181 ( .A1(n7366), .B1(n4639), .ZN(\vrf/N104 ) );
  INR2D0BWP U7182 ( .A1(n7367), .B1(n4639), .ZN(\vrf/N103 ) );
  INR2D0BWP U7183 ( .A1(n7368), .B1(n4639), .ZN(\vrf/N102 ) );
  INR2D0BWP U7184 ( .A1(n7369), .B1(n4643), .ZN(\vrf/N101 ) );
  INR2D0BWP U7185 ( .A1(n7370), .B1(n4631), .ZN(\vrf/N100 ) );
  CKND0BWP U7186 ( .I(n5535), .ZN(n5524) );
  NR4D0BWP U7187 ( .A1(n5544), .A2(n5545), .A3(n5546), .A4(Reset), .ZN(n5535)
         );
  OAI22D0BWP U7188 ( .A1(n5525), .A2(n5541), .B1(n5527), .B2(n5547), .ZN(
        \vrf/N10 ) );
  CKND0BWP U7189 ( .I(instrIn[7]), .ZN(n5547) );
  NR3D0BWP U7190 ( .A1(n5548), .A2(n5549), .A3(n5550), .ZN(n5527) );
  OAI21D0BWP U7191 ( .A1(\srf/N15 ), .A2(n5530), .B(n7436), .ZN(\srf/N59 ) );
  CKND2D0BWP U7192 ( .A1(n5551), .A2(n7438), .ZN(n5530) );
  OAI21D0BWP U7193 ( .A1(\srf/N15 ), .A2(n5532), .B(n7436), .ZN(\srf/N57 ) );
  CKND2D0BWP U7194 ( .A1(\srf/N16 ), .A2(n7438), .ZN(n5532) );
  OAI21D0BWP U7195 ( .A1(\srf/N15 ), .A2(n5533), .B(n7436), .ZN(\srf/N55 ) );
  CKND2D0BWP U7196 ( .A1(\srf/N17 ), .A2(n5551), .ZN(n5533) );
  CKND0BWP U7197 ( .I(\srf/N16 ), .ZN(n5551) );
  OAI21D0BWP U7198 ( .A1(\srf/N15 ), .A2(n5534), .B(n7436), .ZN(\srf/N53 ) );
  AO22D0BWP U7199 ( .A1(scalarWrData[15]), .A2(n5552), .B1(\srf/N20 ), .B2(
        n5553), .Z(\srf/N52 ) );
  AO22D0BWP U7200 ( .A1(scalarWrData[14]), .A2(n5552), .B1(\srf/N21 ), .B2(
        n5553), .Z(\srf/N51 ) );
  AO22D0BWP U7201 ( .A1(scalarWrData[13]), .A2(n5552), .B1(\srf/N22 ), .B2(
        n5553), .Z(\srf/N50 ) );
  AO22D0BWP U7202 ( .A1(scalarWrData[12]), .A2(n5552), .B1(\srf/N23 ), .B2(
        n5553), .Z(\srf/N49 ) );
  AO22D0BWP U7203 ( .A1(scalarWrData[11]), .A2(n5552), .B1(\srf/N24 ), .B2(
        n5553), .Z(\srf/N48 ) );
  AO22D0BWP U7204 ( .A1(scalarWrData[10]), .A2(n5552), .B1(\srf/N25 ), .B2(
        n5553), .Z(\srf/N47 ) );
  AO22D0BWP U7205 ( .A1(scalarWrData[9]), .A2(n5552), .B1(\srf/N26 ), .B2(
        n5553), .Z(\srf/N46 ) );
  AO22D0BWP U7206 ( .A1(scalarWrData[8]), .A2(n5552), .B1(\srf/N27 ), .B2(
        n5553), .Z(\srf/N45 ) );
  AO22D0BWP U7207 ( .A1(scalarWrData[7]), .A2(n5552), .B1(\srf/N28 ), .B2(
        n5553), .Z(\srf/N44 ) );
  AO22D0BWP U7208 ( .A1(scalarWrData[6]), .A2(n5552), .B1(\srf/N29 ), .B2(
        n5553), .Z(\srf/N43 ) );
  AO22D0BWP U7209 ( .A1(scalarWrData[5]), .A2(n5552), .B1(\srf/N30 ), .B2(
        n5553), .Z(\srf/N42 ) );
  AO22D0BWP U7210 ( .A1(scalarWrData[4]), .A2(n5552), .B1(\srf/N31 ), .B2(
        n5553), .Z(\srf/N41 ) );
  AO22D0BWP U7211 ( .A1(scalarWrData[3]), .A2(n5552), .B1(\srf/N32 ), .B2(
        n5553), .Z(\srf/N40 ) );
  AO22D0BWP U7212 ( .A1(scalarWrData[2]), .A2(n5552), .B1(\srf/N33 ), .B2(
        n5553), .Z(\srf/N39 ) );
  AO22D0BWP U7213 ( .A1(scalarWrData[1]), .A2(n5552), .B1(\srf/N34 ), .B2(
        n5553), .Z(\srf/N38 ) );
  AO22D0BWP U7214 ( .A1(scalarWrData[0]), .A2(n5552), .B1(\srf/N35 ), .B2(
        n5553), .Z(\srf/N37 ) );
  NR2D0BWP U7215 ( .A1(n5554), .A2(Reset), .ZN(n5553) );
  NR2D0BWP U7216 ( .A1(n1461), .A2(Reset), .ZN(n5552) );
  CKND2D0BWP U7217 ( .A1(\srf/N16 ), .A2(\srf/N17 ), .ZN(n5534) );
  CKND0BWP U7218 ( .I(\srf/N17 ), .ZN(n7438) );
  CKND0BWP U7219 ( .I(n5555), .ZN(n7439) );
  CKND0BWP U7220 ( .I(n5556), .ZN(n7441) );
  MUX2ND0BWP U7221 ( .I0(n5557), .I1(n5558), .S(N1280), .ZN(n7450) );
  MUX2ND0BWP U7222 ( .I0(n5558), .I1(n5559), .S(N1280), .ZN(n7451) );
  CKND0BWP U7223 ( .I(N1258), .ZN(n5558) );
  MUX2ND0BWP U7224 ( .I0(n5559), .I1(n5560), .S(N1280), .ZN(n7452) );
  CKND0BWP U7225 ( .I(N1259), .ZN(n5559) );
  MUX2ND0BWP U7226 ( .I0(n5560), .I1(n5561), .S(N1280), .ZN(n7453) );
  CKND0BWP U7227 ( .I(N1260), .ZN(n5560) );
  CKND0BWP U7228 ( .I(n5562), .ZN(n7457) );
  CKND0BWP U7229 ( .I(n5563), .ZN(n7458) );
  CKND0BWP U7230 ( .I(n5564), .ZN(n7459) );
  MUX2ND0BWP U7231 ( .I0(n5565), .I1(n5566), .S(\alu/N307 ), .ZN(n7470) );
  MUX2ND0BWP U7232 ( .I0(n5566), .I1(n5567), .S(\alu/N307 ), .ZN(n7471) );
  CKND0BWP U7233 ( .I(\alu/N285 ), .ZN(n5566) );
  MUX2ND0BWP U7234 ( .I0(n5567), .I1(n5568), .S(\alu/N307 ), .ZN(n7472) );
  CKND0BWP U7235 ( .I(\alu/N286 ), .ZN(n5567) );
  MUX2ND0BWP U7236 ( .I0(n5568), .I1(n5569), .S(\alu/N307 ), .ZN(n7473) );
  CKND0BWP U7237 ( .I(\alu/N287 ), .ZN(n5568) );
  CKND0BWP U7238 ( .I(n5570), .ZN(n7475) );
  AOI31D0BWP U7239 ( .A1(n5571), .A2(n5572), .A3(n5573), .B(n5574), .ZN(
        dataOut[9]) );
  NR4D0BWP U7240 ( .A1(n5575), .A2(n5576), .A3(n5577), .A4(n5578), .ZN(n5573)
         );
  OAI22D0BWP U7241 ( .A1(n5579), .A2(n3528), .B1(n5580), .B2(n5581), .ZN(n5578) );
  CKND0BWP U7242 ( .I(vectorData2[105]), .ZN(n5581) );
  OAI22D0BWP U7243 ( .A1(n5582), .A2(n5583), .B1(n5584), .B2(n5585), .ZN(n5577) );
  CKND0BWP U7244 ( .I(vectorData2[73]), .ZN(n5585) );
  CKND0BWP U7245 ( .I(vectorData2[89]), .ZN(n5583) );
  OAI22D0BWP U7246 ( .A1(n5586), .A2(n5587), .B1(n5588), .B2(n5589), .ZN(n5576) );
  CKND0BWP U7247 ( .I(vectorData2[41]), .ZN(n5589) );
  CKND0BWP U7248 ( .I(vectorData2[57]), .ZN(n5587) );
  OAI222D0BWP U7249 ( .A1(n5590), .A2(n3696), .B1(n5591), .B2(n3669), .C1(
        n5592), .C2(n3582), .ZN(n5575) );
  AOI221D0BWP U7250 ( .A1(vectorData2[153]), .A2(n5593), .B1(vectorData2[137]), 
        .B2(n5594), .C(n5595), .ZN(n5572) );
  OAI22D0BWP U7251 ( .A1(n5596), .A2(n3480), .B1(n5597), .B2(n5598), .ZN(n5595) );
  CKND0BWP U7252 ( .I(vectorData2[169]), .ZN(n5598) );
  AOI221D0BWP U7253 ( .A1(vectorData2[233]), .A2(n5599), .B1(vectorData2[249]), 
        .B2(n5600), .C(n5601), .ZN(n5571) );
  OAI22D0BWP U7254 ( .A1(n5602), .A2(n5603), .B1(n5604), .B2(n5605), .ZN(n5601) );
  CKND0BWP U7255 ( .I(vectorData2[217]), .ZN(n5605) );
  CKND0BWP U7256 ( .I(vectorData2[201]), .ZN(n5603) );
  AOI31D0BWP U7257 ( .A1(n5606), .A2(n5607), .A3(n5608), .B(n5574), .ZN(
        dataOut[8]) );
  NR4D0BWP U7258 ( .A1(n5609), .A2(n5610), .A3(n5611), .A4(n5612), .ZN(n5608)
         );
  OAI22D0BWP U7259 ( .A1(n5579), .A2(n3525), .B1(n5580), .B2(n5613), .ZN(n5612) );
  CKND0BWP U7260 ( .I(vectorData2[104]), .ZN(n5613) );
  OAI22D0BWP U7261 ( .A1(n5582), .A2(n5614), .B1(n5584), .B2(n5615), .ZN(n5611) );
  CKND0BWP U7262 ( .I(vectorData2[72]), .ZN(n5615) );
  CKND0BWP U7263 ( .I(vectorData2[88]), .ZN(n5614) );
  OAI22D0BWP U7264 ( .A1(n5586), .A2(n5616), .B1(n5588), .B2(n5617), .ZN(n5610) );
  CKND0BWP U7265 ( .I(vectorData2[40]), .ZN(n5617) );
  CKND0BWP U7266 ( .I(vectorData2[56]), .ZN(n5616) );
  OAI222D0BWP U7267 ( .A1(n5590), .A2(n3693), .B1(n5591), .B2(n3666), .C1(
        n5592), .C2(n3579), .ZN(n5609) );
  AOI221D0BWP U7268 ( .A1(vectorData2[152]), .A2(n5593), .B1(vectorData2[136]), 
        .B2(n5594), .C(n5618), .ZN(n5607) );
  OAI22D0BWP U7269 ( .A1(n5596), .A2(n3477), .B1(n5597), .B2(n5619), .ZN(n5618) );
  CKND0BWP U7270 ( .I(vectorData2[168]), .ZN(n5619) );
  AOI221D0BWP U7271 ( .A1(vectorData2[232]), .A2(n5599), .B1(vectorData2[248]), 
        .B2(n5600), .C(n5620), .ZN(n5606) );
  OAI22D0BWP U7272 ( .A1(n5602), .A2(n5621), .B1(n5604), .B2(n5622), .ZN(n5620) );
  CKND0BWP U7273 ( .I(vectorData2[216]), .ZN(n5622) );
  CKND0BWP U7274 ( .I(vectorData2[200]), .ZN(n5621) );
  AOI31D0BWP U7275 ( .A1(n5623), .A2(n5624), .A3(n5625), .B(n5574), .ZN(
        dataOut[7]) );
  NR4D0BWP U7276 ( .A1(n5626), .A2(n5627), .A3(n5628), .A4(n5629), .ZN(n5625)
         );
  OAI22D0BWP U7277 ( .A1(n5579), .A2(n3558), .B1(n5580), .B2(n5630), .ZN(n5629) );
  CKND0BWP U7278 ( .I(vectorData2[103]), .ZN(n5630) );
  OAI22D0BWP U7279 ( .A1(n5582), .A2(n5631), .B1(n5584), .B2(n5632), .ZN(n5628) );
  CKND0BWP U7280 ( .I(vectorData2[71]), .ZN(n5632) );
  CKND0BWP U7281 ( .I(vectorData2[87]), .ZN(n5631) );
  OAI22D0BWP U7282 ( .A1(n5586), .A2(n5633), .B1(n5588), .B2(n5634), .ZN(n5627) );
  CKND0BWP U7283 ( .I(vectorData2[39]), .ZN(n5634) );
  CKND0BWP U7284 ( .I(vectorData2[55]), .ZN(n5633) );
  OAI222D0BWP U7285 ( .A1(n5590), .A2(n3690), .B1(n5591), .B2(n3663), .C1(
        n5592), .C2(n3612), .ZN(n5626) );
  AOI221D0BWP U7286 ( .A1(vectorData2[151]), .A2(n5593), .B1(vectorData2[135]), 
        .B2(n5594), .C(n5635), .ZN(n5624) );
  OAI22D0BWP U7287 ( .A1(n5596), .A2(n3510), .B1(n5597), .B2(n5636), .ZN(n5635) );
  CKND0BWP U7288 ( .I(vectorData2[167]), .ZN(n5636) );
  AOI221D0BWP U7289 ( .A1(vectorData2[231]), .A2(n5599), .B1(vectorData2[247]), 
        .B2(n5600), .C(n5637), .ZN(n5623) );
  OAI22D0BWP U7290 ( .A1(n5602), .A2(n5638), .B1(n5604), .B2(n5639), .ZN(n5637) );
  CKND0BWP U7291 ( .I(vectorData2[215]), .ZN(n5639) );
  CKND0BWP U7292 ( .I(vectorData2[199]), .ZN(n5638) );
  AOI31D0BWP U7293 ( .A1(n5640), .A2(n5641), .A3(n5642), .B(n5574), .ZN(
        dataOut[6]) );
  NR4D0BWP U7294 ( .A1(n5643), .A2(n5644), .A3(n5645), .A4(n5646), .ZN(n5642)
         );
  OAI22D0BWP U7295 ( .A1(n5579), .A2(n3555), .B1(n5580), .B2(n5647), .ZN(n5646) );
  CKND0BWP U7296 ( .I(vectorData2[102]), .ZN(n5647) );
  OAI22D0BWP U7297 ( .A1(n5582), .A2(n5648), .B1(n5584), .B2(n5649), .ZN(n5645) );
  CKND0BWP U7298 ( .I(vectorData2[70]), .ZN(n5649) );
  CKND0BWP U7299 ( .I(vectorData2[86]), .ZN(n5648) );
  OAI22D0BWP U7300 ( .A1(n5586), .A2(n5650), .B1(n5588), .B2(n5651), .ZN(n5644) );
  CKND0BWP U7301 ( .I(vectorData2[38]), .ZN(n5651) );
  CKND0BWP U7302 ( .I(vectorData2[54]), .ZN(n5650) );
  OAI222D0BWP U7303 ( .A1(n5590), .A2(n3687), .B1(n5591), .B2(n3660), .C1(
        n5592), .C2(n3609), .ZN(n5643) );
  AOI221D0BWP U7304 ( .A1(vectorData2[150]), .A2(n5593), .B1(vectorData2[134]), 
        .B2(n5594), .C(n5652), .ZN(n5641) );
  OAI22D0BWP U7305 ( .A1(n5596), .A2(n3507), .B1(n5597), .B2(n5653), .ZN(n5652) );
  CKND0BWP U7306 ( .I(vectorData2[166]), .ZN(n5653) );
  AOI221D0BWP U7307 ( .A1(vectorData2[230]), .A2(n5599), .B1(vectorData2[246]), 
        .B2(n5600), .C(n5654), .ZN(n5640) );
  OAI22D0BWP U7308 ( .A1(n5602), .A2(n5655), .B1(n5604), .B2(n5656), .ZN(n5654) );
  CKND0BWP U7309 ( .I(vectorData2[214]), .ZN(n5656) );
  CKND0BWP U7310 ( .I(vectorData2[198]), .ZN(n5655) );
  AOI31D0BWP U7311 ( .A1(n5657), .A2(n5658), .A3(n5659), .B(n5574), .ZN(
        dataOut[5]) );
  NR4D0BWP U7312 ( .A1(n5660), .A2(n5661), .A3(n5662), .A4(n5663), .ZN(n5659)
         );
  OAI22D0BWP U7313 ( .A1(n5579), .A2(n3552), .B1(n5580), .B2(n5664), .ZN(n5663) );
  CKND0BWP U7314 ( .I(vectorData2[101]), .ZN(n5664) );
  OAI22D0BWP U7315 ( .A1(n5582), .A2(n5665), .B1(n5584), .B2(n5666), .ZN(n5662) );
  CKND0BWP U7316 ( .I(vectorData2[69]), .ZN(n5666) );
  CKND0BWP U7317 ( .I(vectorData2[85]), .ZN(n5665) );
  OAI22D0BWP U7318 ( .A1(n5586), .A2(n5667), .B1(n5588), .B2(n5668), .ZN(n5661) );
  CKND0BWP U7319 ( .I(vectorData2[37]), .ZN(n5668) );
  CKND0BWP U7320 ( .I(vectorData2[53]), .ZN(n5667) );
  OAI222D0BWP U7321 ( .A1(n5590), .A2(n3684), .B1(n5591), .B2(n3657), .C1(
        n5592), .C2(n3606), .ZN(n5660) );
  AOI221D0BWP U7322 ( .A1(vectorData2[149]), .A2(n5593), .B1(vectorData2[133]), 
        .B2(n5594), .C(n5669), .ZN(n5658) );
  OAI22D0BWP U7323 ( .A1(n5596), .A2(n3504), .B1(n5597), .B2(n5670), .ZN(n5669) );
  CKND0BWP U7324 ( .I(vectorData2[165]), .ZN(n5670) );
  AOI221D0BWP U7325 ( .A1(vectorData2[229]), .A2(n5599), .B1(vectorData2[245]), 
        .B2(n5600), .C(n5671), .ZN(n5657) );
  OAI22D0BWP U7326 ( .A1(n5602), .A2(n5672), .B1(n5604), .B2(n5673), .ZN(n5671) );
  CKND0BWP U7327 ( .I(vectorData2[213]), .ZN(n5673) );
  CKND0BWP U7328 ( .I(vectorData2[197]), .ZN(n5672) );
  AOI31D0BWP U7329 ( .A1(n5674), .A2(n5675), .A3(n5676), .B(n5574), .ZN(
        dataOut[4]) );
  NR4D0BWP U7330 ( .A1(n5677), .A2(n5678), .A3(n5679), .A4(n5680), .ZN(n5676)
         );
  OAI22D0BWP U7331 ( .A1(n5579), .A2(n5681), .B1(n5580), .B2(n3618), .ZN(n5680) );
  CKND0BWP U7332 ( .I(vectorData2[116]), .ZN(n5681) );
  OAI22D0BWP U7333 ( .A1(n5582), .A2(n3516), .B1(n5584), .B2(n3624), .ZN(n5679) );
  OAI22D0BWP U7334 ( .A1(n5586), .A2(n3570), .B1(n5588), .B2(n3462), .ZN(n5678) );
  OAI222D0BWP U7335 ( .A1(n5590), .A2(n5682), .B1(n5591), .B2(n5683), .C1(
        n5592), .C2(n5684), .ZN(n5677) );
  CKND0BWP U7336 ( .I(vectorData2[20]), .ZN(n5684) );
  CKND0BWP U7337 ( .I(vectorData2[4]), .ZN(n5683) );
  CKND0BWP U7338 ( .I(scalarData2[4]), .ZN(n5682) );
  AOI221D0BWP U7339 ( .A1(vectorData2[148]), .A2(n5593), .B1(vectorData2[132]), 
        .B2(n5594), .C(n5685), .ZN(n5675) );
  MOAI22D0BWP U7340 ( .A1(n5597), .A2(n3630), .B1(n5686), .B2(vectorData2[180]), .ZN(n5685) );
  AOI221D0BWP U7341 ( .A1(vectorData2[228]), .A2(n5599), .B1(vectorData2[244]), 
        .B2(n5600), .C(n5687), .ZN(n5674) );
  OAI22D0BWP U7342 ( .A1(n5602), .A2(n3468), .B1(n5604), .B2(n3564), .ZN(n5687) );
  AOI31D0BWP U7343 ( .A1(n5688), .A2(n5689), .A3(n5690), .B(n5574), .ZN(
        dataOut[3]) );
  NR4D0BWP U7344 ( .A1(n5691), .A2(n5692), .A3(n5693), .A4(n5694), .ZN(n5690)
         );
  OAI22D0BWP U7345 ( .A1(n5579), .A2(n5695), .B1(n5580), .B2(n3615), .ZN(n5694) );
  CKND0BWP U7346 ( .I(vectorData2[115]), .ZN(n5695) );
  OAI22D0BWP U7347 ( .A1(n5582), .A2(n3513), .B1(n5584), .B2(n3621), .ZN(n5693) );
  OAI22D0BWP U7348 ( .A1(n5586), .A2(n3567), .B1(n5588), .B2(n3459), .ZN(n5692) );
  OAI222D0BWP U7349 ( .A1(n5590), .A2(n5696), .B1(n5591), .B2(n5697), .C1(
        n5592), .C2(n5698), .ZN(n5691) );
  CKND0BWP U7350 ( .I(vectorData2[19]), .ZN(n5698) );
  CKND0BWP U7351 ( .I(vectorData2[3]), .ZN(n5697) );
  CKND0BWP U7352 ( .I(scalarData2[3]), .ZN(n5696) );
  AOI221D0BWP U7353 ( .A1(vectorData2[147]), .A2(n5593), .B1(vectorData2[131]), 
        .B2(n5594), .C(n5699), .ZN(n5689) );
  MOAI22D0BWP U7354 ( .A1(n5597), .A2(n3627), .B1(n5686), .B2(vectorData2[179]), .ZN(n5699) );
  CKND0BWP U7355 ( .I(n5596), .ZN(n5686) );
  AOI221D0BWP U7356 ( .A1(vectorData2[227]), .A2(n5599), .B1(vectorData2[243]), 
        .B2(n5600), .C(n5700), .ZN(n5688) );
  OAI22D0BWP U7357 ( .A1(n5602), .A2(n3465), .B1(n5604), .B2(n3561), .ZN(n5700) );
  AOI31D0BWP U7358 ( .A1(n5701), .A2(n5702), .A3(n5703), .B(n5574), .ZN(
        dataOut[2]) );
  NR4D0BWP U7359 ( .A1(n5704), .A2(n5705), .A3(n5706), .A4(n5707), .ZN(n5703)
         );
  OAI22D0BWP U7360 ( .A1(n5579), .A2(n3549), .B1(n5580), .B2(n5708), .ZN(n5707) );
  CKND0BWP U7361 ( .I(vectorData2[98]), .ZN(n5708) );
  OAI22D0BWP U7362 ( .A1(n5582), .A2(n5709), .B1(n5584), .B2(n5710), .ZN(n5706) );
  CKND0BWP U7363 ( .I(vectorData2[66]), .ZN(n5710) );
  CKND0BWP U7364 ( .I(vectorData2[82]), .ZN(n5709) );
  OAI22D0BWP U7365 ( .A1(n5586), .A2(n5711), .B1(n5588), .B2(n5712), .ZN(n5705) );
  CKND0BWP U7366 ( .I(vectorData2[34]), .ZN(n5712) );
  CKND0BWP U7367 ( .I(vectorData2[50]), .ZN(n5711) );
  OAI222D0BWP U7368 ( .A1(n5590), .A2(n3681), .B1(n5591), .B2(n3654), .C1(
        n5592), .C2(n3603), .ZN(n5704) );
  AOI221D0BWP U7369 ( .A1(vectorData2[146]), .A2(n5593), .B1(vectorData2[130]), 
        .B2(n5594), .C(n5713), .ZN(n5702) );
  OAI22D0BWP U7370 ( .A1(n5596), .A2(n3501), .B1(n5597), .B2(n5714), .ZN(n5713) );
  CKND0BWP U7371 ( .I(vectorData2[162]), .ZN(n5714) );
  AOI221D0BWP U7372 ( .A1(vectorData2[226]), .A2(n5599), .B1(vectorData2[242]), 
        .B2(n5600), .C(n5715), .ZN(n5701) );
  OAI22D0BWP U7373 ( .A1(n5602), .A2(n5716), .B1(n5604), .B2(n5717), .ZN(n5715) );
  CKND0BWP U7374 ( .I(vectorData2[210]), .ZN(n5717) );
  CKND0BWP U7375 ( .I(vectorData2[194]), .ZN(n5716) );
  AOI31D0BWP U7376 ( .A1(n5718), .A2(n5719), .A3(n5720), .B(n5574), .ZN(
        dataOut[1]) );
  NR4D0BWP U7377 ( .A1(n5721), .A2(n5722), .A3(n5723), .A4(n5724), .ZN(n5720)
         );
  OAI22D0BWP U7378 ( .A1(n5579), .A2(n3522), .B1(n5580), .B2(n5725), .ZN(n5724) );
  CKND0BWP U7379 ( .I(vectorData2[97]), .ZN(n5725) );
  OAI22D0BWP U7380 ( .A1(n5582), .A2(n5726), .B1(n5584), .B2(n5727), .ZN(n5723) );
  CKND0BWP U7381 ( .I(vectorData2[65]), .ZN(n5727) );
  CKND0BWP U7382 ( .I(vectorData2[81]), .ZN(n5726) );
  OAI22D0BWP U7383 ( .A1(n5586), .A2(n5728), .B1(n5588), .B2(n5729), .ZN(n5722) );
  CKND0BWP U7384 ( .I(vectorData2[33]), .ZN(n5729) );
  CKND0BWP U7385 ( .I(vectorData2[49]), .ZN(n5728) );
  OAI222D0BWP U7386 ( .A1(n5590), .A2(n3678), .B1(n5591), .B2(n3651), .C1(
        n5592), .C2(n3576), .ZN(n5721) );
  AOI221D0BWP U7387 ( .A1(vectorData2[145]), .A2(n5593), .B1(vectorData2[129]), 
        .B2(n5594), .C(n5730), .ZN(n5719) );
  OAI22D0BWP U7388 ( .A1(n5596), .A2(n3474), .B1(n5597), .B2(n5731), .ZN(n5730) );
  CKND0BWP U7389 ( .I(vectorData2[161]), .ZN(n5731) );
  AOI221D0BWP U7390 ( .A1(vectorData2[225]), .A2(n5599), .B1(vectorData2[241]), 
        .B2(n5600), .C(n5732), .ZN(n5718) );
  OAI22D0BWP U7391 ( .A1(n5602), .A2(n5733), .B1(n5604), .B2(n5734), .ZN(n5732) );
  CKND0BWP U7392 ( .I(vectorData2[209]), .ZN(n5734) );
  CKND0BWP U7393 ( .I(vectorData2[193]), .ZN(n5733) );
  AOI31D0BWP U7394 ( .A1(n5735), .A2(n5736), .A3(n5737), .B(n5574), .ZN(
        dataOut[15]) );
  NR4D0BWP U7395 ( .A1(n5738), .A2(n5739), .A3(n5740), .A4(n5741), .ZN(n5737)
         );
  OAI22D0BWP U7396 ( .A1(n5579), .A2(n3546), .B1(n5580), .B2(n5742), .ZN(n5741) );
  CKND0BWP U7397 ( .I(vectorData2[111]), .ZN(n5742) );
  OAI22D0BWP U7398 ( .A1(n5582), .A2(n5743), .B1(n5584), .B2(n5744), .ZN(n5740) );
  CKND0BWP U7399 ( .I(vectorData2[79]), .ZN(n5744) );
  CKND0BWP U7400 ( .I(vectorData2[95]), .ZN(n5743) );
  OAI22D0BWP U7401 ( .A1(n5586), .A2(n5745), .B1(n5588), .B2(n5746), .ZN(n5739) );
  CKND0BWP U7402 ( .I(vectorData2[47]), .ZN(n5746) );
  CKND0BWP U7403 ( .I(vectorData2[63]), .ZN(n5745) );
  OAI222D0BWP U7404 ( .A1(n5590), .A2(n5747), .B1(n5591), .B2(n3645), .C1(
        n5592), .C2(n3600), .ZN(n5738) );
  CKND0BWP U7405 ( .I(scalarData2[15]), .ZN(n5747) );
  AOI221D0BWP U7406 ( .A1(vectorData2[159]), .A2(n5593), .B1(vectorData2[143]), 
        .B2(n5594), .C(n5748), .ZN(n5736) );
  OAI22D0BWP U7407 ( .A1(n5596), .A2(n3498), .B1(n5597), .B2(n5749), .ZN(n5748) );
  CKND0BWP U7408 ( .I(vectorData2[175]), .ZN(n5749) );
  AOI221D0BWP U7409 ( .A1(vectorData2[239]), .A2(n5599), .B1(vectorData2[255]), 
        .B2(n5600), .C(n5750), .ZN(n5735) );
  OAI22D0BWP U7410 ( .A1(n5602), .A2(n5751), .B1(n5604), .B2(n5752), .ZN(n5750) );
  CKND0BWP U7411 ( .I(vectorData2[223]), .ZN(n5752) );
  CKND0BWP U7412 ( .I(vectorData2[207]), .ZN(n5751) );
  AOI31D0BWP U7413 ( .A1(n5753), .A2(n5754), .A3(n5755), .B(n5574), .ZN(
        dataOut[14]) );
  NR4D0BWP U7414 ( .A1(n5756), .A2(n5757), .A3(n5758), .A4(n5759), .ZN(n5755)
         );
  OAI22D0BWP U7415 ( .A1(n5579), .A2(n3543), .B1(n5580), .B2(n5760), .ZN(n5759) );
  CKND0BWP U7416 ( .I(vectorData2[110]), .ZN(n5760) );
  OAI22D0BWP U7417 ( .A1(n5582), .A2(n5761), .B1(n5584), .B2(n5762), .ZN(n5758) );
  CKND0BWP U7418 ( .I(vectorData2[78]), .ZN(n5762) );
  CKND0BWP U7419 ( .I(vectorData2[94]), .ZN(n5761) );
  OAI22D0BWP U7420 ( .A1(n5586), .A2(n5763), .B1(n5588), .B2(n5764), .ZN(n5757) );
  CKND0BWP U7421 ( .I(vectorData2[46]), .ZN(n5764) );
  CKND0BWP U7422 ( .I(vectorData2[62]), .ZN(n5763) );
  OAI222D0BWP U7423 ( .A1(n5590), .A2(n5765), .B1(n5591), .B2(n3642), .C1(
        n5592), .C2(n3597), .ZN(n5756) );
  CKND0BWP U7424 ( .I(scalarData2[14]), .ZN(n5765) );
  AOI221D0BWP U7425 ( .A1(vectorData2[158]), .A2(n5593), .B1(vectorData2[142]), 
        .B2(n5594), .C(n5766), .ZN(n5754) );
  OAI22D0BWP U7426 ( .A1(n5596), .A2(n3495), .B1(n5597), .B2(n5767), .ZN(n5766) );
  CKND0BWP U7427 ( .I(vectorData2[174]), .ZN(n5767) );
  AOI221D0BWP U7428 ( .A1(vectorData2[238]), .A2(n5599), .B1(vectorData2[254]), 
        .B2(n5600), .C(n5768), .ZN(n5753) );
  OAI22D0BWP U7429 ( .A1(n5602), .A2(n5769), .B1(n5604), .B2(n5770), .ZN(n5768) );
  CKND0BWP U7430 ( .I(vectorData2[222]), .ZN(n5770) );
  CKND0BWP U7431 ( .I(vectorData2[206]), .ZN(n5769) );
  AOI31D0BWP U7432 ( .A1(n5771), .A2(n5772), .A3(n5773), .B(n5574), .ZN(
        dataOut[13]) );
  NR4D0BWP U7433 ( .A1(n5774), .A2(n5775), .A3(n5776), .A4(n5777), .ZN(n5773)
         );
  OAI22D0BWP U7434 ( .A1(n5579), .A2(n3540), .B1(n5580), .B2(n5778), .ZN(n5777) );
  CKND0BWP U7435 ( .I(vectorData2[109]), .ZN(n5778) );
  OAI22D0BWP U7436 ( .A1(n5582), .A2(n5779), .B1(n5584), .B2(n5780), .ZN(n5776) );
  CKND0BWP U7437 ( .I(vectorData2[77]), .ZN(n5780) );
  CKND0BWP U7438 ( .I(vectorData2[93]), .ZN(n5779) );
  OAI22D0BWP U7439 ( .A1(n5586), .A2(n5781), .B1(n5588), .B2(n5782), .ZN(n5775) );
  CKND0BWP U7440 ( .I(vectorData2[45]), .ZN(n5782) );
  CKND0BWP U7441 ( .I(vectorData2[61]), .ZN(n5781) );
  OAI222D0BWP U7442 ( .A1(n5590), .A2(n5783), .B1(n5591), .B2(n3639), .C1(
        n5592), .C2(n3594), .ZN(n5774) );
  CKND0BWP U7443 ( .I(scalarData2[13]), .ZN(n5783) );
  AOI221D0BWP U7444 ( .A1(vectorData2[157]), .A2(n5593), .B1(vectorData2[141]), 
        .B2(n5594), .C(n5784), .ZN(n5772) );
  OAI22D0BWP U7445 ( .A1(n5596), .A2(n3492), .B1(n5597), .B2(n5785), .ZN(n5784) );
  CKND0BWP U7446 ( .I(vectorData2[173]), .ZN(n5785) );
  AOI221D0BWP U7447 ( .A1(vectorData2[237]), .A2(n5599), .B1(vectorData2[253]), 
        .B2(n5600), .C(n5786), .ZN(n5771) );
  OAI22D0BWP U7448 ( .A1(n5602), .A2(n5787), .B1(n5604), .B2(n5788), .ZN(n5786) );
  CKND0BWP U7449 ( .I(vectorData2[221]), .ZN(n5788) );
  CKND0BWP U7450 ( .I(vectorData2[205]), .ZN(n5787) );
  AOI31D0BWP U7451 ( .A1(n5789), .A2(n5790), .A3(n5791), .B(n5574), .ZN(
        dataOut[12]) );
  NR4D0BWP U7452 ( .A1(n5792), .A2(n5793), .A3(n5794), .A4(n5795), .ZN(n5791)
         );
  OAI22D0BWP U7453 ( .A1(n5579), .A2(n3537), .B1(n5580), .B2(n5796), .ZN(n5795) );
  CKND0BWP U7454 ( .I(vectorData2[108]), .ZN(n5796) );
  OAI22D0BWP U7455 ( .A1(n5582), .A2(n5797), .B1(n5584), .B2(n5798), .ZN(n5794) );
  CKND0BWP U7456 ( .I(vectorData2[76]), .ZN(n5798) );
  CKND0BWP U7457 ( .I(vectorData2[92]), .ZN(n5797) );
  OAI22D0BWP U7458 ( .A1(n5586), .A2(n5799), .B1(n5588), .B2(n5800), .ZN(n5793) );
  CKND0BWP U7459 ( .I(vectorData2[44]), .ZN(n5800) );
  CKND0BWP U7460 ( .I(vectorData2[60]), .ZN(n5799) );
  OAI222D0BWP U7461 ( .A1(n5590), .A2(n5801), .B1(n5591), .B2(n3636), .C1(
        n5592), .C2(n3591), .ZN(n5792) );
  CKND0BWP U7462 ( .I(scalarData2[12]), .ZN(n5801) );
  AOI221D0BWP U7463 ( .A1(vectorData2[156]), .A2(n5593), .B1(vectorData2[140]), 
        .B2(n5594), .C(n5802), .ZN(n5790) );
  OAI22D0BWP U7464 ( .A1(n5596), .A2(n3489), .B1(n5597), .B2(n5803), .ZN(n5802) );
  CKND0BWP U7465 ( .I(vectorData2[172]), .ZN(n5803) );
  AOI221D0BWP U7466 ( .A1(vectorData2[236]), .A2(n5599), .B1(vectorData2[252]), 
        .B2(n5600), .C(n5804), .ZN(n5789) );
  OAI22D0BWP U7467 ( .A1(n5602), .A2(n5805), .B1(n5604), .B2(n5806), .ZN(n5804) );
  CKND0BWP U7468 ( .I(vectorData2[220]), .ZN(n5806) );
  CKND0BWP U7469 ( .I(vectorData2[204]), .ZN(n5805) );
  AOI31D0BWP U7470 ( .A1(n5807), .A2(n5808), .A3(n5809), .B(n5574), .ZN(
        dataOut[11]) );
  NR4D0BWP U7471 ( .A1(n5810), .A2(n5811), .A3(n5812), .A4(n5813), .ZN(n5809)
         );
  OAI22D0BWP U7472 ( .A1(n5579), .A2(n3534), .B1(n5580), .B2(n5814), .ZN(n5813) );
  CKND0BWP U7473 ( .I(vectorData2[107]), .ZN(n5814) );
  OAI22D0BWP U7474 ( .A1(n5582), .A2(n5815), .B1(n5584), .B2(n5816), .ZN(n5812) );
  CKND0BWP U7475 ( .I(vectorData2[75]), .ZN(n5816) );
  CKND0BWP U7476 ( .I(vectorData2[91]), .ZN(n5815) );
  OAI22D0BWP U7477 ( .A1(n5586), .A2(n5817), .B1(n5588), .B2(n5818), .ZN(n5811) );
  CKND0BWP U7478 ( .I(vectorData2[43]), .ZN(n5818) );
  CKND0BWP U7479 ( .I(vectorData2[59]), .ZN(n5817) );
  OAI222D0BWP U7480 ( .A1(n5590), .A2(n5819), .B1(n5591), .B2(n3633), .C1(
        n5592), .C2(n3588), .ZN(n5810) );
  CKND0BWP U7481 ( .I(scalarData2[11]), .ZN(n5819) );
  AOI221D0BWP U7482 ( .A1(vectorData2[155]), .A2(n5593), .B1(vectorData2[139]), 
        .B2(n5594), .C(n5820), .ZN(n5808) );
  OAI22D0BWP U7483 ( .A1(n5596), .A2(n3486), .B1(n5597), .B2(n5821), .ZN(n5820) );
  CKND0BWP U7484 ( .I(vectorData2[171]), .ZN(n5821) );
  AOI221D0BWP U7485 ( .A1(vectorData2[235]), .A2(n5599), .B1(vectorData2[251]), 
        .B2(n5600), .C(n5822), .ZN(n5807) );
  OAI22D0BWP U7486 ( .A1(n5602), .A2(n5823), .B1(n5604), .B2(n5824), .ZN(n5822) );
  CKND0BWP U7487 ( .I(vectorData2[219]), .ZN(n5824) );
  CKND0BWP U7488 ( .I(vectorData2[203]), .ZN(n5823) );
  AOI31D0BWP U7489 ( .A1(n5825), .A2(n5826), .A3(n5827), .B(n5574), .ZN(
        dataOut[10]) );
  NR4D0BWP U7490 ( .A1(n5828), .A2(n5829), .A3(n5830), .A4(n5831), .ZN(n5827)
         );
  OAI22D0BWP U7491 ( .A1(n5579), .A2(n3531), .B1(n5580), .B2(n5832), .ZN(n5831) );
  CKND0BWP U7492 ( .I(vectorData2[106]), .ZN(n5832) );
  OAI22D0BWP U7493 ( .A1(n5582), .A2(n5833), .B1(n5584), .B2(n5834), .ZN(n5830) );
  CKND0BWP U7494 ( .I(vectorData2[74]), .ZN(n5834) );
  CKND0BWP U7495 ( .I(vectorData2[90]), .ZN(n5833) );
  OAI22D0BWP U7496 ( .A1(n5586), .A2(n5835), .B1(n5588), .B2(n5836), .ZN(n5829) );
  CKND0BWP U7497 ( .I(vectorData2[42]), .ZN(n5836) );
  CKND0BWP U7498 ( .I(vectorData2[58]), .ZN(n5835) );
  OAI222D0BWP U7499 ( .A1(n5590), .A2(n3699), .B1(n5591), .B2(n3672), .C1(
        n5592), .C2(n3585), .ZN(n5828) );
  AOI221D0BWP U7500 ( .A1(vectorData2[154]), .A2(n5593), .B1(vectorData2[138]), 
        .B2(n5594), .C(n5837), .ZN(n5826) );
  OAI22D0BWP U7501 ( .A1(n5596), .A2(n3483), .B1(n5597), .B2(n5838), .ZN(n5837) );
  CKND0BWP U7502 ( .I(vectorData2[170]), .ZN(n5838) );
  AOI221D0BWP U7503 ( .A1(vectorData2[234]), .A2(n5599), .B1(vectorData2[250]), 
        .B2(n5600), .C(n5839), .ZN(n5825) );
  OAI22D0BWP U7504 ( .A1(n5602), .A2(n5840), .B1(n5604), .B2(n5841), .ZN(n5839) );
  CKND0BWP U7505 ( .I(vectorData2[218]), .ZN(n5841) );
  CKND0BWP U7506 ( .I(vectorData2[202]), .ZN(n5840) );
  AOI31D0BWP U7507 ( .A1(n5842), .A2(n5843), .A3(n5844), .B(n5574), .ZN(
        dataOut[0]) );
  NR4D0BWP U7508 ( .A1(n5845), .A2(n5846), .A3(n5847), .A4(n5848), .ZN(n5844)
         );
  OAI22D0BWP U7509 ( .A1(n5579), .A2(n3519), .B1(n5580), .B2(n5849), .ZN(n5848) );
  CKND0BWP U7510 ( .I(vectorData2[96]), .ZN(n5849) );
  OAI22D0BWP U7511 ( .A1(n5582), .A2(n5850), .B1(n5584), .B2(n5851), .ZN(n5847) );
  CKND0BWP U7512 ( .I(vectorData2[64]), .ZN(n5851) );
  CKND0BWP U7513 ( .I(vectorData2[80]), .ZN(n5850) );
  OAI22D0BWP U7514 ( .A1(n5586), .A2(n5852), .B1(n5588), .B2(n5853), .ZN(n5846) );
  CKND0BWP U7515 ( .I(vectorData2[32]), .ZN(n5853) );
  CKND0BWP U7516 ( .I(vectorData2[48]), .ZN(n5852) );
  OAI222D0BWP U7517 ( .A1(n5590), .A2(n3675), .B1(n5591), .B2(n3648), .C1(
        n5592), .C2(n3573), .ZN(n5845) );
  ND3D0BWP U7518 ( .A1(n5592), .A2(n5854), .A3(n5855), .ZN(n5591) );
  ND3D0BWP U7519 ( .A1(n5855), .A2(n5592), .A3(n5548), .ZN(n5590) );
  CKND0BWP U7520 ( .I(n5854), .ZN(n5548) );
  CKND2D0BWP U7521 ( .A1(n5856), .A2(n5857), .ZN(n5592) );
  AN4D0BWP U7522 ( .A1(n5858), .A2(n5588), .A3(n5859), .A4(n5860), .Z(n5855)
         );
  NR4D0BWP U7523 ( .A1(n5861), .A2(n5594), .A3(n5600), .A4(n5599), .ZN(n5860)
         );
  ND4D0BWP U7524 ( .A1(n5604), .A2(n5602), .A3(n5597), .A4(n5862), .ZN(n5861)
         );
  AN4D0BWP U7525 ( .A1(n5596), .A2(n5579), .A3(n5580), .A4(n5582), .Z(n5859)
         );
  ND3D0BWP U7526 ( .A1(n5856), .A2(n5863), .A3(cycles[2]), .ZN(n5582) );
  CKND2D0BWP U7527 ( .A1(n5864), .A2(cycles[1]), .ZN(n5580) );
  CKND2D0BWP U7528 ( .A1(n5865), .A2(n5863), .ZN(n5579) );
  ND3D0BWP U7529 ( .A1(n5857), .A2(n5866), .A3(cycles[1]), .ZN(n5588) );
  AN2D0BWP U7530 ( .A1(n5584), .A2(n5586), .Z(n5858) );
  CKND2D0BWP U7531 ( .A1(n5867), .A2(n5857), .ZN(n5586) );
  CKND2D0BWP U7532 ( .A1(n5864), .A2(n5868), .ZN(n5584) );
  INR3D0BWP U7533 ( .A1(n5863), .B1(cycles[0]), .B2(n5869), .ZN(n5864) );
  AOI221D0BWP U7534 ( .A1(vectorData2[144]), .A2(n5593), .B1(vectorData2[128]), 
        .B2(n5594), .C(n5870), .ZN(n5843) );
  OAI22D0BWP U7535 ( .A1(n5596), .A2(n3471), .B1(n5597), .B2(n5871), .ZN(n5870) );
  CKND0BWP U7536 ( .I(vectorData2[160]), .ZN(n5871) );
  ND3D0BWP U7537 ( .A1(n5872), .A2(n5869), .A3(cycles[1]), .ZN(n5597) );
  CKND0BWP U7538 ( .I(n5874), .ZN(n5867) );
  INR3D0BWP U7539 ( .A1(n5872), .B1(cycles[1]), .B2(cycles[2]), .ZN(n5594) );
  CKND0BWP U7540 ( .I(n5862), .ZN(n5593) );
  ND4D0BWP U7541 ( .A1(cycles[3]), .A2(n5856), .A3(n5869), .A4(n5873), .ZN(
        n5862) );
  AOI221D0BWP U7542 ( .A1(vectorData2[224]), .A2(n5599), .B1(vectorData2[240]), 
        .B2(n5600), .C(n5875), .ZN(n5842) );
  OAI22D0BWP U7543 ( .A1(n5602), .A2(n5876), .B1(n5604), .B2(n5877), .ZN(n5875) );
  CKND0BWP U7544 ( .I(vectorData2[208]), .ZN(n5877) );
  IND3D0BWP U7545 ( .A1(n5878), .B1(n5873), .B2(n5856), .ZN(n5604) );
  CKND0BWP U7546 ( .I(vectorData2[192]), .ZN(n5876) );
  ND3D0BWP U7547 ( .A1(n5872), .A2(n5868), .A3(cycles[2]), .ZN(n5602) );
  INR3D0BWP U7548 ( .A1(n5872), .B1(n5868), .B2(n5869), .ZN(n5599) );
  NR3D0BWP U7549 ( .A1(cycles[0]), .A2(cycles[4]), .A3(n5879), .ZN(n5872) );
  CKND2D0BWP U7550 ( .A1(n5880), .A2(n5881), .ZN(\alu/N999 ) );
  OAI22D0BWP U7551 ( .A1(n5882), .A2(n5883), .B1(n5884), .B2(n5885), .ZN(
        \alu/N991 ) );
  CKND0BWP U7552 ( .I(\alu/N849 ), .ZN(n5884) );
  OAI22D0BWP U7553 ( .A1(n5883), .A2(n5885), .B1(n5882), .B2(n5886), .ZN(
        \alu/N990 ) );
  CKND0BWP U7554 ( .I(\alu/N848 ), .ZN(n5883) );
  OAI22D0BWP U7555 ( .A1(n5885), .A2(n5886), .B1(n5882), .B2(n5887), .ZN(
        \alu/N989 ) );
  CKND0BWP U7556 ( .I(\alu/N847 ), .ZN(n5886) );
  OAI22D0BWP U7557 ( .A1(n5885), .A2(n5887), .B1(n5882), .B2(n5888), .ZN(
        \alu/N988 ) );
  CKND0BWP U7558 ( .I(\alu/N846 ), .ZN(n5887) );
  OAI22D0BWP U7559 ( .A1(n5885), .A2(n5888), .B1(n5882), .B2(n5889), .ZN(
        \alu/N987 ) );
  CKND0BWP U7560 ( .I(\alu/N845 ), .ZN(n5888) );
  OAI22D0BWP U7561 ( .A1(n5885), .A2(n5889), .B1(n5882), .B2(n5890), .ZN(
        \alu/N986 ) );
  CKND0BWP U7562 ( .I(\alu/N844 ), .ZN(n5889) );
  OAI22D0BWP U7563 ( .A1(n5885), .A2(n5890), .B1(n5882), .B2(n5891), .ZN(
        \alu/N985 ) );
  CKND0BWP U7564 ( .I(\alu/N843 ), .ZN(n5890) );
  OAI22D0BWP U7565 ( .A1(n5885), .A2(n5891), .B1(n5882), .B2(n5892), .ZN(
        \alu/N984 ) );
  CKND0BWP U7566 ( .I(\alu/N842 ), .ZN(n5891) );
  OAI22D0BWP U7567 ( .A1(n5885), .A2(n5892), .B1(n5882), .B2(n5893), .ZN(
        \alu/N983 ) );
  CKND0BWP U7568 ( .I(n5894), .ZN(n5882) );
  CKND0BWP U7569 ( .I(\alu/N841 ), .ZN(n5892) );
  MOAI22D0BWP U7570 ( .A1(n5885), .A2(n5893), .B1(\alu/N839 ), .B2(n5894), 
        .ZN(\alu/N982 ) );
  NR2D0BWP U7571 ( .A1(\alu/N850 ), .A2(n5895), .ZN(n5894) );
  CKND0BWP U7572 ( .I(\alu/N840 ), .ZN(n5893) );
  CKND2D0BWP U7573 ( .A1(n5880), .A2(n5896), .ZN(\alu/N836 ) );
  CKND2D0BWP U7574 ( .A1(n5880), .A2(n5897), .ZN(\alu/N835 ) );
  CKND2D0BWP U7575 ( .A1(n5880), .A2(n5898), .ZN(\alu/N834 ) );
  CKND2D0BWP U7576 ( .A1(n5880), .A2(n5899), .ZN(\alu/N833 ) );
  CKND0BWP U7577 ( .I(\alu/N997 ), .ZN(n5880) );
  INR2D0BWP U7578 ( .A1(\U3/U27/Z_0 ), .B1(n5895), .ZN(\alu/N814 ) );
  OAI221D0BWP U7579 ( .A1(n5900), .A2(n5896), .B1(n5901), .B2(n5902), .C(n5903), .ZN(\alu/N665 ) );
  OAI221D0BWP U7580 ( .A1(n5904), .A2(n5902), .B1(n5900), .B2(n5897), .C(n5903), .ZN(\alu/N664 ) );
  OAI221D0BWP U7581 ( .A1(n5905), .A2(n5902), .B1(n5900), .B2(n5898), .C(n5903), .ZN(\alu/N663 ) );
  OAI221D0BWP U7582 ( .A1(n5906), .A2(n5902), .B1(n5900), .B2(n5899), .C(n5903), .ZN(\alu/N662 ) );
  CKND0BWP U7583 ( .I(\alu/N540 ), .ZN(n5899) );
  OAI221D0BWP U7584 ( .A1(n5900), .A2(n5881), .B1(n5902), .B2(n5907), .C(n5903), .ZN(\alu/N661 ) );
  CKND0BWP U7585 ( .I(n5908), .ZN(n5903) );
  CKND0BWP U7586 ( .I(n5909), .ZN(n5907) );
  CKND0BWP U7587 ( .I(n5910), .ZN(n5902) );
  CKND0BWP U7588 ( .I(\alu/N539 ), .ZN(n5881) );
  NR2D0BWP U7589 ( .A1(n5911), .A2(n5912), .ZN(n5900) );
  NR2D0BWP U7590 ( .A1(n5913), .A2(n5908), .ZN(\alu/N660 ) );
  AOI222D0BWP U7591 ( .A1(n5914), .A2(n5912), .B1(n7460), .B2(n5910), .C1(
        \alu/N610 ), .C2(n5911), .ZN(n5913) );
  NR2D0BWP U7592 ( .A1(n5915), .A2(n5908), .ZN(\alu/N659 ) );
  AOI222D0BWP U7593 ( .A1(n7460), .A2(n5912), .B1(n5910), .B2(\alu/N529 ), 
        .C1(\alu/N609 ), .C2(n5911), .ZN(n5915) );
  NR2D0BWP U7594 ( .A1(n5916), .A2(n5908), .ZN(\alu/N658 ) );
  AOI222D0BWP U7595 ( .A1(n5912), .A2(\alu/N529 ), .B1(n7467), .B2(n5910), 
        .C1(\alu/N608 ), .C2(n5911), .ZN(n5916) );
  NR2D0BWP U7596 ( .A1(n5917), .A2(n5908), .ZN(\alu/N657 ) );
  AOI222D0BWP U7597 ( .A1(n7467), .A2(n5912), .B1(n7466), .B2(n5910), .C1(
        \alu/N607 ), .C2(n5911), .ZN(n5917) );
  NR2D0BWP U7598 ( .A1(n5918), .A2(n5908), .ZN(\alu/N656 ) );
  AOI222D0BWP U7599 ( .A1(n7466), .A2(n5912), .B1(n7465), .B2(n5910), .C1(
        \alu/N606 ), .C2(n5911), .ZN(n5918) );
  NR2D0BWP U7600 ( .A1(n5919), .A2(n5908), .ZN(\alu/N655 ) );
  AOI222D0BWP U7601 ( .A1(n7465), .A2(n5912), .B1(n7464), .B2(n5910), .C1(
        \alu/N605 ), .C2(n5911), .ZN(n5919) );
  NR2D0BWP U7602 ( .A1(n5920), .A2(n5908), .ZN(\alu/N654 ) );
  AOI222D0BWP U7603 ( .A1(n7464), .A2(n5912), .B1(n7463), .B2(n5910), .C1(
        \alu/N604 ), .C2(n5911), .ZN(n5920) );
  NR2D0BWP U7604 ( .A1(n5921), .A2(n5908), .ZN(\alu/N653 ) );
  AOI222D0BWP U7605 ( .A1(n7463), .A2(n5912), .B1(n7462), .B2(n5910), .C1(
        \alu/N603 ), .C2(n5911), .ZN(n5921) );
  NR2D0BWP U7606 ( .A1(n5922), .A2(n5908), .ZN(\alu/N652 ) );
  AOI222D0BWP U7607 ( .A1(n7462), .A2(n5912), .B1(n7461), .B2(n5910), .C1(
        \alu/N602 ), .C2(n5911), .ZN(n5922) );
  NR2D0BWP U7608 ( .A1(n5923), .A2(n5908), .ZN(\alu/N651 ) );
  ND4D0BWP U7609 ( .A1(n5924), .A2(n5925), .A3(n5926), .A4(n5927), .ZN(n5908)
         );
  INR2D0BWP U7610 ( .A1(n5928), .B1(n5929), .ZN(n5926) );
  ND4D0BWP U7611 ( .A1(n5930), .A2(n5931), .A3(n5932), .A4(n5933), .ZN(n5925)
         );
  INR3D0BWP U7612 ( .A1(n5934), .B1(n5935), .B2(n5936), .ZN(n5933) );
  MUX2ND0BWP U7613 ( .I0(n5937), .I1(n5938), .S(n5939), .ZN(n5932) );
  CKND2D0BWP U7614 ( .A1(n5940), .A2(n5941), .ZN(n5938) );
  CKND2D0BWP U7615 ( .A1(n5942), .A2(n5943), .ZN(n5937) );
  ND4D0BWP U7616 ( .A1(\alu/N539 ), .A2(n5912), .A3(\alu/N540 ), .A4(n5944), 
        .ZN(n5924) );
  NR3D0BWP U7617 ( .A1(n5896), .A2(n5898), .A3(n5897), .ZN(n5944) );
  CKND0BWP U7618 ( .I(\alu/N542 ), .ZN(n5897) );
  CKND0BWP U7619 ( .I(\alu/N541 ), .ZN(n5898) );
  CKND0BWP U7620 ( .I(\alu/N543 ), .ZN(n5896) );
  AOI222D0BWP U7621 ( .A1(n7461), .A2(n5912), .B1(n5910), .B2(\alu/N521 ), 
        .C1(\alu/N601 ), .C2(n5911), .ZN(n5923) );
  NR2D0BWP U7622 ( .A1(n5945), .A2(n5912), .ZN(n5910) );
  CKMUX2D0BWP U7623 ( .I0(op1[15]), .I1(op2[15]), .S(n5946), .Z(\alu/N634 ) );
  INR2D0BWP U7624 ( .A1(n5927), .B1(n5947), .ZN(n5946) );
  CKND0BWP U7625 ( .I(n5935), .ZN(n7468) );
  MUX2ND0BWP U7626 ( .I0(n5949), .I1(n5950), .S(\alu/N307 ), .ZN(\alu/N443 )
         );
  MUX2ND0BWP U7627 ( .I0(n5951), .I1(n5949), .S(\alu/N307 ), .ZN(\alu/N442 )
         );
  CKND0BWP U7628 ( .I(\alu/N293 ), .ZN(n5949) );
  MUX2ND0BWP U7629 ( .I0(n5952), .I1(n5951), .S(\alu/N307 ), .ZN(\alu/N441 )
         );
  CKND0BWP U7630 ( .I(\alu/N292 ), .ZN(n5951) );
  MUX2ND0BWP U7631 ( .I0(n5953), .I1(n5952), .S(\alu/N307 ), .ZN(\alu/N440 )
         );
  CKND0BWP U7632 ( .I(\alu/N291 ), .ZN(n5952) );
  MUX2ND0BWP U7633 ( .I0(n5954), .I1(n5953), .S(\alu/N307 ), .ZN(\alu/N439 )
         );
  CKND0BWP U7634 ( .I(\alu/N290 ), .ZN(n5953) );
  MUX2ND0BWP U7635 ( .I0(n5569), .I1(n5954), .S(\alu/N307 ), .ZN(\alu/N438 )
         );
  CKND0BWP U7636 ( .I(\alu/N289 ), .ZN(n5954) );
  CKND0BWP U7637 ( .I(\alu/N288 ), .ZN(n5569) );
  MUX2ND0BWP U7638 ( .I0(n5955), .I1(n5565), .S(\alu/N307 ), .ZN(\alu/N433 )
         );
  CKND0BWP U7639 ( .I(\alu/N284 ), .ZN(n5565) );
  MUX2ND0BWP U7640 ( .I0(n5956), .I1(n5955), .S(\alu/N307 ), .ZN(\alu/N432 )
         );
  CKND0BWP U7641 ( .I(\alu/N283 ), .ZN(n5955) );
  MUX2ND0BWP U7642 ( .I0(n5957), .I1(n5956), .S(\alu/N307 ), .ZN(\alu/N431 )
         );
  CKND0BWP U7643 ( .I(\alu/N282 ), .ZN(n5956) );
  CKND0BWP U7644 ( .I(n5958), .ZN(\alu/N376 ) );
  CKND0BWP U7645 ( .I(n5959), .ZN(\alu/N311 ) );
  CKND0BWP U7646 ( .I(n5960), .ZN(\alu/N310 ) );
  CKND0BWP U7647 ( .I(n5961), .ZN(\alu/N309 ) );
  CKND0BWP U7648 ( .I(n5962), .ZN(\alu/N308 ) );
  CKXOR2D0BWP U7649 ( .A1(n5963), .A2(\U3/U27/Z_0 ), .Z(\alu/N1019 ) );
  XOR3D0BWP U7650 ( .A1(op2[14]), .A2(n5964), .A3(n5965), .Z(\alu/N1018 ) );
  XOR3D0BWP U7651 ( .A1(op2[13]), .A2(n5966), .A3(n5967), .Z(\alu/N1017 ) );
  XOR3D0BWP U7652 ( .A1(op2[12]), .A2(n5968), .A3(n5969), .Z(\alu/N1016 ) );
  XOR3D0BWP U7653 ( .A1(op2[11]), .A2(n5970), .A3(n5971), .Z(\alu/N1015 ) );
  XOR3D0BWP U7654 ( .A1(op2[10]), .A2(n5972), .A3(n5973), .Z(\alu/N1014 ) );
  XOR3D0BWP U7655 ( .A1(op2[9]), .A2(n5974), .A3(n5975), .Z(\alu/N1013 ) );
  XOR3D0BWP U7656 ( .A1(op2[8]), .A2(n5976), .A3(n5977), .Z(\alu/N1012 ) );
  XOR3D0BWP U7657 ( .A1(op2[7]), .A2(n5978), .A3(n3370), .Z(\alu/N1011 ) );
  XOR3D0BWP U7658 ( .A1(op2[6]), .A2(op1[6]), .A3(n5979), .Z(\alu/N1010 ) );
  XOR3D0BWP U7659 ( .A1(op2[5]), .A2(op1[5]), .A3(n5980), .Z(\alu/N1009 ) );
  XOR3D0BWP U7660 ( .A1(op2[4]), .A2(op1[4]), .A3(n5981), .Z(\alu/N1008 ) );
  XOR3D0BWP U7661 ( .A1(op2[3]), .A2(op1[3]), .A3(n5982), .Z(\alu/N1007 ) );
  XOR3D0BWP U7662 ( .A1(op2[2]), .A2(op1[2]), .A3(n5983), .Z(\alu/N1006 ) );
  XNR3D0BWP U7663 ( .A1(op2[1]), .A2(op1[1]), .A3(n5984), .ZN(\alu/N1005 ) );
  CKND2D0BWP U7664 ( .A1(op2[0]), .A2(op1[0]), .ZN(n5984) );
  CKXOR2D0BWP U7665 ( .A1(op2[0]), .A2(op1[0]), .Z(\alu/N1004 ) );
  NR2D0BWP U7666 ( .A1(n5985), .A2(n5539), .ZN(addrDst[2]) );
  CKND0BWP U7667 ( .I(instrIn[11]), .ZN(n5539) );
  NR2D0BWP U7668 ( .A1(n5985), .A2(n5541), .ZN(addrDst[1]) );
  CKND0BWP U7669 ( .I(instrIn[10]), .ZN(n5541) );
  NR2D0BWP U7670 ( .A1(n5985), .A2(n5526), .ZN(addrDst[0]) );
  CKND0BWP U7671 ( .I(instrIn[9]), .ZN(n5526) );
  AN3D0BWP U7672 ( .A1(n5546), .A2(n5986), .A3(n5525), .Z(n5985) );
  CKXOR2D0BWP U7673 ( .A1(scalarToLoad[15]), .A2(result[15]), .Z(\U3/U8/Z_0 )
         );
  CKMUX2D0BWP U7674 ( .I0(N1168), .I1(N1169), .S(n5988), .Z(\U3/U6/Z_25 ) );
  MUX2ND0BWP U7675 ( .I0(n5989), .I1(n3390), .S(n5987), .ZN(\U3/U6/Z_24 ) );
  MUX2ND0BWP U7676 ( .I0(n5990), .I1(n3391), .S(n5987), .ZN(\U3/U6/Z_23 ) );
  MUX2ND0BWP U7677 ( .I0(n5991), .I1(n3382), .S(n5987), .ZN(\U3/U6/Z_22 ) );
  MUX2ND0BWP U7678 ( .I0(n5992), .I1(n3383), .S(n5987), .ZN(\U3/U6/Z_21 ) );
  MUX2ND0BWP U7679 ( .I0(n5993), .I1(n3384), .S(n5987), .ZN(\U3/U6/Z_20 ) );
  MUX2ND0BWP U7680 ( .I0(n5994), .I1(n3385), .S(n5987), .ZN(\U3/U6/Z_19 ) );
  MUX2ND0BWP U7681 ( .I0(n5995), .I1(n3386), .S(n5987), .ZN(\U3/U6/Z_18 ) );
  MUX2ND0BWP U7682 ( .I0(n5996), .I1(n3387), .S(n5987), .ZN(\U3/U6/Z_17 ) );
  MUX2ND0BWP U7683 ( .I0(n5997), .I1(n3388), .S(n5987), .ZN(\U3/U6/Z_16 ) );
  MUX2ND0BWP U7684 ( .I0(n5998), .I1(n3389), .S(n5987), .ZN(\U3/U6/Z_15 ) );
  OAI211D0BWP U7685 ( .A1(n5999), .A2(n6000), .B(n6001), .C(n6002), .ZN(
        \U3/U32/Z_0 ) );
  CKND2D0BWP U7686 ( .A1(n5947), .A2(n6003), .ZN(n6000) );
  NR3D0BWP U7687 ( .A1(n5999), .A2(n5947), .A3(n5885), .ZN(\U3/U31/Z_0 ) );
  CKND2D0BWP U7688 ( .A1(\alu/N850 ), .A2(n6003), .ZN(n5885) );
  OAI22D0BWP U7689 ( .A1(n6004), .A2(n6005), .B1(n5928), .B2(n6006), .ZN(
        \U3/U30/Z_4 ) );
  OAI21D0BWP U7690 ( .A1(n5967), .A2(n6007), .B(n6008), .ZN(\U3/U30/Z_3 ) );
  MUX2ND0BWP U7691 ( .I0(n6009), .I1(n6010), .S(op2[13]), .ZN(n6008) );
  OAI21D0BWP U7692 ( .A1(n6011), .A2(n6006), .B(n6004), .ZN(n6010) );
  INR2D0BWP U7693 ( .A1(n6011), .B1(n6006), .ZN(n6009) );
  OAI21D0BWP U7694 ( .A1(n5969), .A2(n6007), .B(n6012), .ZN(\U3/U30/Z_2 ) );
  MUX2ND0BWP U7695 ( .I0(n6013), .I1(n6014), .S(op2[12]), .ZN(n6012) );
  AO21D0BWP U7696 ( .A1(n6015), .A2(n6016), .B(n6017), .Z(n6014) );
  NR3D0BWP U7697 ( .A1(n6006), .A2(n6018), .A3(n6015), .ZN(n6013) );
  OAI21D0BWP U7698 ( .A1(n5971), .A2(n6007), .B(n6019), .ZN(\U3/U30/Z_1 ) );
  MUX2ND0BWP U7699 ( .I0(n6020), .I1(n6017), .S(op2[11]), .ZN(n6019) );
  OAI21D0BWP U7700 ( .A1(op2[10]), .A2(n6006), .B(n6004), .ZN(n6017) );
  CKND0BWP U7701 ( .I(n6021), .ZN(n6004) );
  NR2D0BWP U7702 ( .A1(n6018), .A2(n6006), .ZN(n6020) );
  CKND0BWP U7703 ( .I(n6016), .ZN(n6006) );
  OAI21D0BWP U7704 ( .A1(n5973), .A2(n6007), .B(n6022), .ZN(\U3/U30/Z_0 ) );
  MUX2ND0BWP U7705 ( .I0(n6016), .I1(n6021), .S(op2[10]), .ZN(n6022) );
  OAI21D0BWP U7706 ( .A1(n6023), .A2(n6024), .B(n6001), .ZN(n6021) );
  NR2D0BWP U7707 ( .A1(n6024), .A2(n5947), .ZN(n6016) );
  OAI32D0BWP U7708 ( .A1(n6025), .A2(n6026), .A3(n6027), .B1(n5965), .B2(n6001), .ZN(\U3/U29/Z_4 ) );
  OAI22D0BWP U7709 ( .A1(n5967), .A2(n6001), .B1(n6026), .B2(n6028), .ZN(
        \U3/U29/Z_3 ) );
  XNR2D0BWP U7710 ( .A1(n6025), .A2(n6027), .ZN(n6028) );
  OA22D1BWP U7711 ( .A1(n5967), .A2(n5999), .B1(n6029), .B2(n6030), .Z(n6027)
         );
  ND3D0BWP U7712 ( .A1(n6031), .A2(n6032), .A3(n6033), .ZN(n6025) );
  OAI22D0BWP U7713 ( .A1(n5969), .A2(n6001), .B1(n6026), .B2(n6034), .ZN(
        \U3/U29/Z_2 ) );
  XNR2D0BWP U7714 ( .A1(n6033), .A2(n6035), .ZN(n6034) );
  AN2D0BWP U7715 ( .A1(n6031), .A2(n6032), .Z(n6035) );
  OAI22D0BWP U7716 ( .A1(n5969), .A2(n5999), .B1(n6029), .B2(n6036), .ZN(n6033) );
  OAI22D0BWP U7717 ( .A1(n5971), .A2(n6001), .B1(n6026), .B2(n6037), .ZN(
        \U3/U29/Z_1 ) );
  XNR2D0BWP U7718 ( .A1(n6032), .A2(n6031), .ZN(n6037) );
  OAI22D0BWP U7719 ( .A1(n5971), .A2(n5999), .B1(n6029), .B2(n6015), .ZN(n6031) );
  OAI22D0BWP U7720 ( .A1(n5973), .A2(n6001), .B1(n6026), .B2(n6032), .ZN(
        \U3/U29/Z_0 ) );
  OAI22D0BWP U7721 ( .A1(n5973), .A2(n5999), .B1(n6029), .B2(n6018), .ZN(n6032) );
  AN2D0BWP U7722 ( .A1(n6038), .A2(n6039), .Z(n6029) );
  CKND2D0BWP U7723 ( .A1(\alu/N851 ), .A2(n6040), .ZN(n5999) );
  AN2D0BWP U7724 ( .A1(n6024), .A2(n6007), .Z(n6026) );
  AO21D0BWP U7725 ( .A1(n6038), .A2(n6039), .B(n5895), .Z(n6007) );
  CKND0BWP U7726 ( .I(n6003), .ZN(n5895) );
  CKND2D0BWP U7727 ( .A1(n6041), .A2(n6042), .ZN(n6039) );
  CKND2D0BWP U7728 ( .A1(n6043), .A2(n6042), .ZN(n6038) );
  CKXOR2D0BWP U7729 ( .A1(op1[15]), .A2(op2[15]), .Z(\U3/U27/Z_0 ) );
  CKND2D0BWP U7730 ( .A1(n6044), .A2(n5947), .ZN(\U3/U25/Z_25 ) );
  MUX2ND0BWP U7731 ( .I0(n6045), .I1(n5975), .S(n5947), .ZN(\U3/U25/Z_24 ) );
  MUX2ND0BWP U7732 ( .I0(n6046), .I1(n5977), .S(n5947), .ZN(\U3/U25/Z_23 ) );
  MUX2ND0BWP U7733 ( .I0(n3374), .I1(n3370), .S(n5947), .ZN(\U3/U25/Z_22 ) );
  MUX2ND0BWP U7734 ( .I0(n3372), .I1(n3380), .S(n5947), .ZN(\U3/U25/Z_21 ) );
  MUX2ND0BWP U7735 ( .I0(n3378), .I1(n3377), .S(n5947), .ZN(\U3/U25/Z_20 ) );
  MUX2ND0BWP U7736 ( .I0(n3373), .I1(n3376), .S(n5947), .ZN(\U3/U25/Z_19 ) );
  MUX2ND0BWP U7737 ( .I0(n3375), .I1(n3381), .S(n5947), .ZN(\U3/U25/Z_18 ) );
  MUX2ND0BWP U7738 ( .I0(n3379), .I1(n3371), .S(n5947), .ZN(\U3/U25/Z_17 ) );
  CKMUX2D0BWP U7739 ( .I0(op1[1]), .I1(op2[1]), .S(n6023), .Z(\U3/U25/Z_16 )
         );
  MUX2ND0BWP U7740 ( .I0(n6047), .I1(n6048), .S(n5947), .ZN(\U3/U25/Z_15 ) );
  OAI21D0BWP U7741 ( .A1(n5563), .A2(n6049), .B(n6050), .ZN(\U3/U23/Z_3 ) );
  ND4D0BWP U7742 ( .A1(n6051), .A2(n6052), .A3(n6053), .A4(n6054), .ZN(n5563)
         );
  CKND2D0BWP U7743 ( .A1(n6055), .A2(n6056), .ZN(n6054) );
  AO21D0BWP U7744 ( .A1(\U3/U24/Z_0 ), .A2(\alu/N579 ), .B(n6040), .Z(
        \U3/U23/Z_2 ) );
  OAI21D0BWP U7745 ( .A1(n6049), .A2(n5564), .B(n6050), .ZN(\U3/U23/Z_1 ) );
  CKND2D0BWP U7746 ( .A1(n6053), .A2(n6057), .ZN(n5564) );
  OAI31D0BWP U7747 ( .A1(n7466), .A2(n6058), .A3(n7465), .B(n6052), .ZN(n6057)
         );
  AOI211D0BWP U7748 ( .A1(n6055), .A2(\alu/N521 ), .B(n7464), .C(n7463), .ZN(
        n6058) );
  AO221D0BWP U7749 ( .A1(n6059), .A2(n5912), .B1(\alu/N600 ), .B2(\U3/U24/Z_0 ), .C(n6040), .Z(\U3/U23/Z_0 ) );
  AOI21D0BWP U7750 ( .A1(n6061), .A2(n6062), .B(n7467), .ZN(n6060) );
  OAI21D0BWP U7751 ( .A1(n6063), .A2(n7464), .B(n6064), .ZN(n6062) );
  AOI21D0BWP U7752 ( .A1(n7461), .A2(n6065), .B(n7463), .ZN(n6063) );
  AO21D0BWP U7753 ( .A1(n214), .A2(n6040), .B(n6066), .Z(\U3/U22/Z_5 ) );
  AO221D0BWP U7754 ( .A1(n6067), .A2(n6068), .B1(n215), .B2(n6040), .C(n6066), 
        .Z(\U3/U22/Z_4 ) );
  CKND0BWP U7755 ( .I(n5901), .ZN(n6067) );
  MUX2ND0BWP U7756 ( .I0(n5942), .I1(n5941), .S(n6069), .ZN(n5901) );
  XNR2D0BWP U7757 ( .A1(n5941), .A2(n6070), .ZN(n5942) );
  CKND2D0BWP U7758 ( .A1(n6071), .A2(n6072), .ZN(n6070) );
  OAI22D0BWP U7759 ( .A1(n6073), .A2(n6074), .B1(n6075), .B2(n6076), .ZN(n5941) );
  CKND0BWP U7760 ( .I(\alu/N312 ), .ZN(n6073) );
  OAI21D0BWP U7761 ( .A1(n6023), .A2(n5965), .B(n6005), .ZN(\alu/N312 ) );
  MOAI22D0BWP U7762 ( .A1(n6077), .A2(n5904), .B1(n216), .B2(n6078), .ZN(
        \U3/U22/Z_3 ) );
  MUX2ND0BWP U7763 ( .I0(n6072), .I1(n5930), .S(n5948), .ZN(n5904) );
  XNR2D0BWP U7764 ( .A1(n6072), .A2(n6079), .ZN(n5930) );
  CKND2D0BWP U7765 ( .A1(n6071), .A2(n5943), .ZN(n6079) );
  OAI22D0BWP U7766 ( .A1(n5959), .A2(n6074), .B1(n6075), .B2(n6080), .ZN(n6072) );
  MUX2ND0BWP U7767 ( .I0(op2[13]), .I1(op1[13]), .S(n5947), .ZN(n5959) );
  MOAI22D0BWP U7768 ( .A1(n6077), .A2(n5905), .B1(n217), .B2(n6078), .ZN(
        \U3/U22/Z_2 ) );
  MUX2ND0BWP U7769 ( .I0(n6081), .I1(n5931), .S(n5948), .ZN(n5905) );
  MAOI22D0BWP U7770 ( .A1(n5943), .A2(n6071), .B1(n6082), .B2(n6081), .ZN(
        n5931) );
  AN2D0BWP U7771 ( .A1(n6083), .A2(n6084), .Z(n6082) );
  AN3D0BWP U7772 ( .A1(n6083), .A2(n5939), .A3(n6081), .Z(n6071) );
  OAI22D0BWP U7773 ( .A1(n5960), .A2(n6074), .B1(n6075), .B2(n6085), .ZN(n6081) );
  MUX2ND0BWP U7774 ( .I0(op2[12]), .I1(op1[12]), .S(n5947), .ZN(n5960) );
  MOAI22D0BWP U7775 ( .A1(n6077), .A2(n5906), .B1(n218), .B2(n6078), .ZN(
        \U3/U22/Z_1 ) );
  CKND2D0BWP U7776 ( .A1(n6024), .A2(n6002), .ZN(n6078) );
  CKND2D0BWP U7777 ( .A1(n6042), .A2(n6086), .ZN(n6002) );
  NR2D0BWP U7778 ( .A1(n5947), .A2(\alu/N851 ), .ZN(n6042) );
  OAI211D0BWP U7779 ( .A1(n6041), .A2(n6043), .B(n6003), .C(\alu/N851 ), .ZN(
        n6024) );
  MUX2ND0BWP U7780 ( .I0(n6083), .I1(n5934), .S(n5948), .ZN(n5906) );
  CKXOR2D0BWP U7781 ( .A1(n6084), .A2(n6083), .Z(n5934) );
  AN2D0BWP U7782 ( .A1(n5939), .A2(n5943), .Z(n6084) );
  OAI22D0BWP U7783 ( .A1(n5961), .A2(n6074), .B1(n6075), .B2(n6087), .ZN(n6083) );
  CKND0BWP U7784 ( .I(\alu/N421 ), .ZN(n6087) );
  MUX2ND0BWP U7785 ( .I0(op2[11]), .I1(op1[11]), .S(n5947), .ZN(n5961) );
  AO221D0BWP U7786 ( .A1(n5909), .A2(n6068), .B1(n219), .B2(n6040), .C(n6066), 
        .Z(\U3/U22/Z_0 ) );
  INR2D0BWP U7787 ( .A1(n6088), .B1(n6050), .ZN(n6066) );
  OAI21D0BWP U7788 ( .A1(\alu/N851 ), .A2(n6023), .B(n6003), .ZN(n6088) );
  CKND0BWP U7789 ( .I(n6077), .ZN(n6068) );
  AOI21D0BWP U7790 ( .A1(n6059), .A2(n5912), .B(\U3/U24/Z_0 ), .ZN(n6077) );
  CKND0BWP U7791 ( .I(n6049), .ZN(\U3/U24/Z_0 ) );
  CKND2D0BWP U7792 ( .A1(n5911), .A2(n6059), .ZN(n6049) );
  INR2D0BWP U7793 ( .A1(n6089), .B1(n5914), .ZN(n5911) );
  CKND0BWP U7794 ( .I(n5945), .ZN(n5914) );
  MUX2ND0BWP U7795 ( .I0(\alu/N456 ), .I1(\alu/N476 ), .S(n5948), .ZN(n5945)
         );
  AO211D0BWP U7796 ( .A1(\alu/N419 ), .A2(n6090), .B(\alu/N338 ), .C(
        \alu/N307 ), .Z(\alu/N456 ) );
  AOI31D0BWP U7797 ( .A1(n6051), .A2(n6052), .A3(n6091), .B(n5912), .ZN(n6089)
         );
  INR3D0BWP U7798 ( .A1(n6055), .B1(n7460), .B2(\alu/N521 ), .ZN(n6091) );
  CKND0BWP U7799 ( .I(n6056), .ZN(\alu/N521 ) );
  MUX2ND0BWP U7800 ( .I0(\alu/N446 ), .I1(\alu/N466 ), .S(n5948), .ZN(n6056)
         );
  CKND0BWP U7801 ( .I(n6053), .ZN(n7460) );
  MUX2ND0BWP U7802 ( .I0(\alu/N455 ), .I1(\alu/N475 ), .S(n5948), .ZN(n6053)
         );
  AO222D0BWP U7803 ( .A1(\alu/N418 ), .A2(n6090), .B1(\alu/N337 ), .B2(n6092), 
        .C1(\alu/N338 ), .C2(\alu/N307 ), .Z(\alu/N455 ) );
  NR2D0BWP U7804 ( .A1(n7462), .A2(n7461), .ZN(n6055) );
  AO222D0BWP U7805 ( .A1(\alu/N410 ), .A2(n6090), .B1(\alu/N329 ), .B2(n6092), 
        .C1(\alu/N330 ), .C2(\alu/N307 ), .Z(\alu/N447 ) );
  CKND0BWP U7806 ( .I(n6065), .ZN(n7462) );
  MUX2ND0BWP U7807 ( .I0(\alu/N448 ), .I1(\alu/N468 ), .S(n5948), .ZN(n6065)
         );
  AO222D0BWP U7808 ( .A1(\alu/N411 ), .A2(n6090), .B1(\alu/N330 ), .B2(n6092), 
        .C1(\alu/N331 ), .C2(\alu/N307 ), .Z(\alu/N448 ) );
  NR2D0BWP U7809 ( .A1(n7467), .A2(\alu/N529 ), .ZN(n6052) );
  AO222D0BWP U7810 ( .A1(\alu/N417 ), .A2(n6090), .B1(\alu/N336 ), .B2(n6092), 
        .C1(\alu/N337 ), .C2(\alu/N307 ), .Z(\alu/N454 ) );
  AO222D0BWP U7811 ( .A1(\alu/N416 ), .A2(n6090), .B1(\alu/N335 ), .B2(n6092), 
        .C1(\alu/N336 ), .C2(\alu/N307 ), .Z(\alu/N453 ) );
  NR4D0BWP U7812 ( .A1(n7466), .A2(n7465), .A3(n7464), .A4(n7463), .ZN(n6051)
         );
  AO222D0BWP U7813 ( .A1(\alu/N412 ), .A2(n6090), .B1(\alu/N331 ), .B2(n6092), 
        .C1(\alu/N332 ), .C2(\alu/N307 ), .Z(\alu/N449 ) );
  AO222D0BWP U7814 ( .A1(\alu/N413 ), .A2(n6090), .B1(\alu/N332 ), .B2(n6092), 
        .C1(\alu/N333 ), .C2(\alu/N307 ), .Z(\alu/N450 ) );
  CKND0BWP U7815 ( .I(n6064), .ZN(n7465) );
  MUX2ND0BWP U7816 ( .I0(\alu/N451 ), .I1(\alu/N471 ), .S(n5948), .ZN(n6064)
         );
  AO222D0BWP U7817 ( .A1(\alu/N414 ), .A2(n6090), .B1(\alu/N333 ), .B2(n6092), 
        .C1(\alu/N334 ), .C2(\alu/N307 ), .Z(\alu/N451 ) );
  CKND0BWP U7818 ( .I(n6061), .ZN(n7466) );
  MUX2ND0BWP U7819 ( .I0(\alu/N452 ), .I1(\alu/N472 ), .S(n5948), .ZN(n6061)
         );
  AO222D0BWP U7820 ( .A1(\alu/N415 ), .A2(n6090), .B1(\alu/N334 ), .B2(n6092), 
        .C1(\alu/N335 ), .C2(\alu/N307 ), .Z(\alu/N452 ) );
  XNR2D0BWP U7821 ( .A1(n5939), .A2(n6069), .ZN(n5909) );
  CKND2D0BWP U7822 ( .A1(n5943), .A2(n5948), .ZN(n6069) );
  AN4D0BWP U7823 ( .A1(n6093), .A2(n6094), .A3(n6095), .A4(n6096), .Z(n5936)
         );
  NR4D0BWP U7824 ( .A1(\alu/N293 ), .A2(\alu/N292 ), .A3(\alu/N291 ), .A4(
        \alu/N290 ), .ZN(n6096) );
  NR4D0BWP U7825 ( .A1(\alu/N289 ), .A2(\alu/N288 ), .A3(\alu/N287 ), .A4(
        \alu/N286 ), .ZN(n6095) );
  NR4D0BWP U7826 ( .A1(\alu/N285 ), .A2(\alu/N284 ), .A3(\alu/N283 ), .A4(
        \alu/N282 ), .ZN(n6094) );
  NR3D0BWP U7827 ( .A1(n6097), .A2(n7469), .A3(\alu/N446 ), .ZN(n6093) );
  AO222D0BWP U7828 ( .A1(\alu/N409 ), .A2(n6090), .B1(\alu/N328 ), .B2(n6092), 
        .C1(\alu/N329 ), .C2(\alu/N307 ), .Z(\alu/N446 ) );
  AO222D0BWP U7829 ( .A1(\alu/N407 ), .A2(n6090), .B1(\alu/N326 ), .B2(n6092), 
        .C1(\alu/N327 ), .C2(\alu/N307 ), .Z(n7469) );
  MUX2ND0BWP U7830 ( .I0(n5957), .I1(n5950), .S(\alu/N307 ), .ZN(n6097) );
  CKND0BWP U7831 ( .I(\alu/N326 ), .ZN(n5950) );
  CKND0BWP U7832 ( .I(\alu/N281 ), .ZN(n5957) );
  AOI222D0BWP U7833 ( .A1(\alu/N328 ), .A2(\alu/N307 ), .B1(\alu/N408 ), .B2(
        n6090), .C1(\alu/N327 ), .C2(n6092), .ZN(n5935) );
  CKND2D0BWP U7834 ( .A1(n6098), .A2(n6074), .ZN(n6092) );
  AN4D0BWP U7835 ( .A1(\alu/N420 ), .A2(\alu/N307 ), .A3(\alu/N421 ), .A4(
        n6099), .Z(n5929) );
  NR3D0BWP U7836 ( .A1(n6076), .A2(n6085), .A3(n6080), .ZN(n6099) );
  CKND0BWP U7837 ( .I(\alu/N423 ), .ZN(n6080) );
  CKND0BWP U7838 ( .I(\alu/N422 ), .ZN(n6085) );
  CKND0BWP U7839 ( .I(\alu/N424 ), .ZN(n6076) );
  CKND0BWP U7840 ( .I(n5940), .ZN(n5943) );
  IIND4D0BWP U7841 ( .A1(\alu/N466 ), .A2(\alu/N467 ), .B1(n6100), .B2(n6101), 
        .ZN(n5940) );
  NR4D0BWP U7842 ( .A1(n6102), .A2(\alu/N473 ), .A3(\alu/N475 ), .A4(
        \alu/N474 ), .ZN(n6101) );
  OR2D0BWP U7843 ( .A1(\alu/N471 ), .A2(\alu/N472 ), .Z(n6102) );
  NR3D0BWP U7844 ( .A1(\alu/N468 ), .A2(\alu/N470 ), .A3(\alu/N469 ), .ZN(
        n6100) );
  OAI22D0BWP U7845 ( .A1(n5962), .A2(n6074), .B1(n6075), .B2(n6103), .ZN(n5939) );
  CKND0BWP U7846 ( .I(\alu/N420 ), .ZN(n6103) );
  NR2D0BWP U7847 ( .A1(n6090), .A2(\alu/N307 ), .ZN(n6075) );
  INR3D0BWP U7848 ( .A1(n6098), .B1(\alu/N307 ), .B2(\alu/N338 ), .ZN(n6090)
         );
  ND4D0BWP U7849 ( .A1(n6104), .A2(n6105), .A3(n6106), .A4(n6107), .ZN(n6098)
         );
  NR2D0BWP U7850 ( .A1(\alu/N337 ), .A2(\alu/N307 ), .ZN(n6106) );
  CKND2D0BWP U7851 ( .A1(\alu/N338 ), .A2(n7474), .ZN(n6074) );
  CKND0BWP U7852 ( .I(\alu/N307 ), .ZN(n7474) );
  MUX2ND0BWP U7853 ( .I0(op2[10]), .I1(op1[10]), .S(n5947), .ZN(n5962) );
  NR2D0BWP U7854 ( .A1(n5965), .A2(n6001), .ZN(n6110) );
  OAI32D0BWP U7855 ( .A1(n6001), .A2(op2[14]), .A3(n5965), .B1(n6111), .B2(
        n6112), .ZN(n6109) );
  MOAI22D0BWP U7856 ( .A1(n6036), .A2(n6113), .B1(op2[13]), .B2(n6114), .ZN(
        n6112) );
  OAI32D0BWP U7857 ( .A1(n6115), .A2(n6116), .A3(n6015), .B1(n6117), .B2(n6118), .ZN(n6111) );
  OAI21D0BWP U7858 ( .A1(n5973), .A2(n6001), .B(n6119), .ZN(n6118) );
  AOI21D0BWP U7859 ( .A1(op2[10]), .A2(n6120), .B(n6011), .ZN(n6117) );
  OAI22D0BWP U7860 ( .A1(n6015), .A2(n6113), .B1(n6116), .B2(n6115), .ZN(n6120) );
  INR2D0BWP U7861 ( .A1(n6113), .B1(op2[12]), .ZN(n6116) );
  OAI21D0BWP U7862 ( .A1(n5969), .A2(n6001), .B(n6119), .ZN(n6113) );
  OAI21D0BWP U7863 ( .A1(n5971), .A2(n6001), .B(n6119), .ZN(n6115) );
  NR2D0BWP U7864 ( .A1(op2[13]), .A2(n6114), .ZN(n6108) );
  AOI21D0BWP U7865 ( .A1(op1[13]), .A2(n6059), .B(n6086), .ZN(n6114) );
  CKND0BWP U7866 ( .I(n6119), .ZN(n6086) );
  CKND2D0BWP U7867 ( .A1(n6003), .A2(n6040), .ZN(n6119) );
  CKND0BWP U7868 ( .I(n6050), .ZN(n6040) );
  NR2D0BWP U7869 ( .A1(n6041), .A2(n6043), .ZN(n6050) );
  AN3D0BWP U7870 ( .A1(n6121), .A2(n5485), .A3(func[0]), .Z(n6043) );
  NR4D0BWP U7871 ( .A1(n6122), .A2(func[0]), .A3(func[2]), .A4(func[3]), .ZN(
        n6041) );
  OAI22D0BWP U7872 ( .A1(n6123), .A2(n6044), .B1(n6124), .B2(n6125), .ZN(n6003) );
  CKND0BWP U7873 ( .I(\alu/N88 ), .ZN(n6125) );
  ND4D0BWP U7874 ( .A1(n6030), .A2(n6005), .A3(n6036), .A4(n6126), .ZN(
        \alu/N88 ) );
  NR2D0BWP U7875 ( .A1(op2[11]), .A2(op2[10]), .ZN(n6126) );
  NR4D0BWP U7876 ( .A1(n6127), .A2(n6128), .A3(op2[1]), .A4(op2[0]), .ZN(n6124) );
  ND3D0BWP U7877 ( .A1(n3375), .A2(n3373), .A3(n3379), .ZN(n6128) );
  ND4D0BWP U7878 ( .A1(n3378), .A2(n3372), .A3(n6129), .A4(n3374), .ZN(n6127)
         );
  NR2D0BWP U7879 ( .A1(op2[9]), .A2(op2[8]), .ZN(n6129) );
  CKND0BWP U7880 ( .I(\alu/N87 ), .ZN(n6044) );
  ND4D0BWP U7881 ( .A1(n5969), .A2(n5967), .A3(n5971), .A4(n6130), .ZN(
        \alu/N87 ) );
  NR2D0BWP U7882 ( .A1(op1[10]), .A2(\alu/N851 ), .ZN(n6130) );
  NR4D0BWP U7883 ( .A1(n6131), .A2(n6132), .A3(op1[1]), .A4(op1[0]), .ZN(n6123) );
  ND3D0BWP U7884 ( .A1(n3381), .A2(n3376), .A3(n3371), .ZN(n6132) );
  ND4D0BWP U7885 ( .A1(n3377), .A2(n3380), .A3(n6133), .A4(n3370), .ZN(n6131)
         );
  NR2D0BWP U7886 ( .A1(op1[9]), .A2(op1[8]), .ZN(n6133) );
  CKND0BWP U7887 ( .I(n6001), .ZN(n6059) );
  ND4D0BWP U7888 ( .A1(n6121), .A2(n5927), .A3(n6134), .A4(n5928), .ZN(n6001)
         );
  ND3D0BWP U7889 ( .A1(op2[14]), .A2(op2[13]), .A3(n6011), .ZN(n5928) );
  NR3D0BWP U7890 ( .A1(n6015), .A2(n6018), .A3(n6036), .ZN(n6011) );
  NR2D0BWP U7891 ( .A1(func[3]), .A2(func[0]), .ZN(n6134) );
  ND4D0BWP U7892 ( .A1(\alu/N851 ), .A2(op1[13]), .A3(n6135), .A4(op1[12]), 
        .ZN(n5927) );
  NR2D0BWP U7893 ( .A1(n5973), .A2(n5971), .ZN(n6135) );
  NR2D0BWP U7894 ( .A1(\alu/N307 ), .A2(n5958), .ZN(\U3/U19/Z_3 ) );
  IND4D0BWP U7895 ( .A1(n6105), .B1(n6104), .B2(n6107), .B3(n6136), .ZN(n5958)
         );
  NR3D0BWP U7896 ( .A1(\alu/N329 ), .A2(\alu/N330 ), .A3(\alu/N328 ), .ZN(
        n6105) );
  INR2D0BWP U7897 ( .A1(\alu/N385 ), .B1(\alu/N307 ), .ZN(\U3/U19/Z_2 ) );
  NR4D0BWP U7898 ( .A1(\alu/N331 ), .A2(\alu/N332 ), .A3(\alu/N333 ), .A4(
        \alu/N334 ), .ZN(n6104) );
  NR2D0BWP U7899 ( .A1(\alu/N307 ), .A2(n5570), .ZN(\U3/U19/Z_1 ) );
  CKND2D0BWP U7900 ( .A1(n6136), .A2(n6137), .ZN(n5570) );
  OAI31D0BWP U7901 ( .A1(n6138), .A2(\alu/N334 ), .A3(\alu/N333 ), .B(n6107), 
        .ZN(n6137) );
  NR2D0BWP U7902 ( .A1(\alu/N335 ), .A2(\alu/N336 ), .ZN(n6107) );
  AOI211D0BWP U7903 ( .A1(n6139), .A2(\alu/N328 ), .B(\alu/N332 ), .C(
        \alu/N331 ), .ZN(n6138) );
  NR2D0BWP U7904 ( .A1(\alu/N330 ), .A2(\alu/N329 ), .ZN(n6139) );
  OR2D0BWP U7905 ( .A1(\alu/N406 ), .A2(\alu/N307 ), .Z(\U3/U19/Z_0 ) );
  CKND0BWP U7906 ( .I(\alu/N337 ), .ZN(n6136) );
  AOI21D0BWP U7907 ( .A1(n6141), .A2(n6142), .B(\alu/N335 ), .ZN(n6140) );
  CKND0BWP U7908 ( .I(\alu/N334 ), .ZN(n6142) );
  OAI21D0BWP U7909 ( .A1(\alu/N332 ), .A2(n6143), .B(n6144), .ZN(n6141) );
  CKND0BWP U7910 ( .I(\alu/N333 ), .ZN(n6144) );
  AOI21D0BWP U7911 ( .A1(\alu/N329 ), .A2(n6145), .B(\alu/N331 ), .ZN(n6143)
         );
  CKND0BWP U7912 ( .I(\alu/N330 ), .ZN(n6145) );
  NR2D0BWP U7913 ( .A1(n6146), .A2(n5555), .ZN(\U3/U17/Z_3 ) );
  OAI31D0BWP U7914 ( .A1(n7442), .A2(n7443), .A3(N1602), .B(n6147), .ZN(n5555)
         );
  INR2D0BWP U7915 ( .A1(N1660), .B1(n6146), .ZN(\U3/U17/Z_2 ) );
  NR2D0BWP U7916 ( .A1(n6146), .A2(n5556), .ZN(\U3/U17/Z_1 ) );
  OAI31D0BWP U7917 ( .A1(n7448), .A2(n6148), .A3(N1610), .B(n6149), .ZN(n5556)
         );
  AOI211D0BWP U7918 ( .A1(n6150), .A2(n6151), .B(n7447), .C(n7446), .ZN(n6148)
         );
  AOI31D0BWP U7919 ( .A1(N1602), .A2(n6152), .A3(n6153), .B(n7444), .ZN(n6150)
         );
  OAI221D0BWP U7920 ( .A1(n6154), .A2(n6155), .B1(n6156), .B2(n6146), .C(n6157), .ZN(\U3/U17/Z_0 ) );
  CKND0BWP U7921 ( .I(N1681), .ZN(n6156) );
  OAI22D0BWP U7922 ( .A1(n6158), .A2(n5873), .B1(n6159), .B2(n6160), .ZN(
        \U3/U16/Z_4 ) );
  OAI22D0BWP U7923 ( .A1(n6158), .A2(n5879), .B1(n6159), .B2(n6161), .ZN(
        \U3/U16/Z_3 ) );
  OAI22D0BWP U7924 ( .A1(n6158), .A2(n5869), .B1(n6159), .B2(n6162), .ZN(
        \U3/U16/Z_2 ) );
  OAI22D0BWP U7925 ( .A1(n6158), .A2(n5868), .B1(n6159), .B2(n6163), .ZN(
        \U3/U16/Z_1 ) );
  OAI22D0BWP U7926 ( .A1(n6158), .A2(n5866), .B1(n6159), .B2(n6164), .ZN(
        \U3/U16/Z_0 ) );
  AOI21D0BWP U7927 ( .A1(n6165), .A2(n6166), .B(n7440), .ZN(n6159) );
  CKND0BWP U7928 ( .I(n6146), .ZN(n7440) );
  CKND2D0BWP U7929 ( .A1(n6167), .A2(n6165), .ZN(n6146) );
  OA21D0BWP U7930 ( .A1(n6168), .A2(n6169), .B(n6170), .Z(n6158) );
  NR2D0BWP U7931 ( .A1(n6171), .A2(n5873), .ZN(\U3/U14/Z_4 ) );
  CKND0BWP U7932 ( .I(cycles[4]), .ZN(n5873) );
  OAI22D0BWP U7933 ( .A1(n6171), .A2(n5879), .B1(n6172), .B2(n6173), .ZN(
        \U3/U14/Z_3 ) );
  MOAI22D0BWP U7934 ( .A1(n6171), .A2(n5869), .B1(n7456), .B2(N1466), .ZN(
        \U3/U14/Z_2 ) );
  OAI22D0BWP U7935 ( .A1(n6171), .A2(n5868), .B1(n6172), .B2(n5562), .ZN(
        \U3/U14/Z_1 ) );
  CKND2D0BWP U7936 ( .A1(n6174), .A2(n6175), .ZN(n5562) );
  OAI31D0BWP U7937 ( .A1(n6176), .A2(N1415), .A3(N1414), .B(n6177), .ZN(n6175)
         );
  AOI211D0BWP U7938 ( .A1(n6178), .A2(N1409), .B(N1413), .C(N1412), .ZN(n6176)
         );
  NR2D0BWP U7939 ( .A1(N1411), .A2(N1410), .ZN(n6178) );
  OAI211D0BWP U7940 ( .A1(n6179), .A2(n6154), .B(n6180), .C(n6181), .ZN(
        \U3/U14/Z_0 ) );
  MAOI22D0BWP U7941 ( .A1(n7456), .A2(N1487), .B1(n5866), .B2(n6171), .ZN(
        n6181) );
  OAI22D0BWP U7942 ( .A1(n6180), .A2(n3398), .B1(n6171), .B2(n5989), .ZN(
        \U3/U13/Z_9 ) );
  OAI22D0BWP U7943 ( .A1(n6180), .A2(n3399), .B1(n6171), .B2(n5990), .ZN(
        \U3/U13/Z_8 ) );
  OAI22D0BWP U7944 ( .A1(n6180), .A2(n3400), .B1(n6171), .B2(n5991), .ZN(
        \U3/U13/Z_7 ) );
  OAI22D0BWP U7945 ( .A1(n6180), .A2(n3401), .B1(n6171), .B2(n5992), .ZN(
        \U3/U13/Z_6 ) );
  OAI22D0BWP U7946 ( .A1(n6180), .A2(n3402), .B1(n6171), .B2(n5993), .ZN(
        \U3/U13/Z_5 ) );
  OAI222D0BWP U7947 ( .A1(n6171), .A2(n5994), .B1(n6182), .B2(n6183), .C1(
        n6180), .C2(n3420), .ZN(\U3/U13/Z_4 ) );
  OAI222D0BWP U7948 ( .A1(n6171), .A2(n5995), .B1(n6182), .B2(n6184), .C1(
        n6180), .C2(n3421), .ZN(\U3/U13/Z_3 ) );
  OAI222D0BWP U7949 ( .A1(n6171), .A2(n5996), .B1(n6182), .B2(n6185), .C1(
        n6180), .C2(n3422), .ZN(\U3/U13/Z_2 ) );
  OAI22D0BWP U7950 ( .A1(n6180), .A2(n3392), .B1(n6171), .B2(n6186), .ZN(
        \U3/U13/Z_15 ) );
  OAI22D0BWP U7951 ( .A1(n6180), .A2(n3393), .B1(n6171), .B2(n6187), .ZN(
        \U3/U13/Z_14 ) );
  OAI22D0BWP U7952 ( .A1(n6180), .A2(n3394), .B1(n6171), .B2(n6188), .ZN(
        \U3/U13/Z_13 ) );
  OAI22D0BWP U7953 ( .A1(n6180), .A2(n3395), .B1(n6171), .B2(n6189), .ZN(
        \U3/U13/Z_12 ) );
  OAI22D0BWP U7954 ( .A1(n6180), .A2(n3396), .B1(n6171), .B2(n6190), .ZN(
        \U3/U13/Z_11 ) );
  OAI22D0BWP U7955 ( .A1(n6180), .A2(n3397), .B1(n6171), .B2(n6191), .ZN(
        \U3/U13/Z_10 ) );
  OAI222D0BWP U7956 ( .A1(n6171), .A2(n5997), .B1(n6182), .B2(n6192), .C1(
        n6180), .C2(n3423), .ZN(\U3/U13/Z_1 ) );
  OAI222D0BWP U7957 ( .A1(n6171), .A2(n5998), .B1(n6182), .B2(n6193), .C1(
        n6180), .C2(n3424), .ZN(\U3/U13/Z_0 ) );
  AOI21D0BWP U7958 ( .A1(N1280), .A2(n6165), .B(n7456), .ZN(n6182) );
  CKND2D0BWP U7959 ( .A1(n6165), .A2(n6194), .ZN(n6172) );
  CKND0BWP U7960 ( .I(n6154), .ZN(n6165) );
  CKND2D0BWP U7961 ( .A1(n6195), .A2(n6196), .ZN(n6154) );
  CKND2D0BWP U7962 ( .A1(n3266), .A2(n6197), .ZN(RD) );
  OAI31D0BWP U7963 ( .A1(n5544), .A2(n5546), .A3(n5545), .B(n1461), .ZN(N4366)
         );
  CKND0BWP U7964 ( .I(n5554), .ZN(n1461) );
  AOI211D0BWP U7965 ( .A1(n5525), .A2(n5986), .B(n5545), .C(n5544), .ZN(n5554)
         );
  AOI21D0BWP U7966 ( .A1(n6198), .A2(n6199), .B(n6200), .ZN(n5546) );
  AO222D0BWP U7967 ( .A1(N572), .A2(n4659), .B1(N2882), .B2(n4693), .C1(n4742), 
        .C2(n7197), .Z(N4364) );
  AO222D0BWP U7968 ( .A1(N571), .A2(n4659), .B1(N2881), .B2(n4693), .C1(n4742), 
        .C2(n7198), .Z(N4363) );
  AO222D0BWP U7969 ( .A1(N570), .A2(n4659), .B1(N2880), .B2(n4693), .C1(n4742), 
        .C2(n7199), .Z(N4362) );
  AO222D0BWP U7970 ( .A1(N569), .A2(n4659), .B1(N2879), .B2(n4693), .C1(n4742), 
        .C2(n7200), .Z(N4361) );
  AO222D0BWP U7971 ( .A1(N568), .A2(n4659), .B1(N2878), .B2(n4693), .C1(n4742), 
        .C2(n7201), .Z(N4360) );
  AO222D0BWP U7972 ( .A1(N567), .A2(n4659), .B1(N2877), .B2(n4693), .C1(n4742), 
        .C2(n7202), .Z(N4359) );
  AO222D0BWP U7973 ( .A1(N566), .A2(n4659), .B1(N2876), .B2(n4693), .C1(n4742), 
        .C2(n7203), .Z(N4358) );
  AO222D0BWP U7974 ( .A1(N565), .A2(n4659), .B1(N2875), .B2(n4693), .C1(n4742), 
        .C2(n7204), .Z(N4357) );
  AO222D0BWP U7975 ( .A1(N564), .A2(n4659), .B1(N2874), .B2(n4693), .C1(n4742), 
        .C2(n7205), .Z(N4356) );
  AO222D0BWP U7976 ( .A1(N563), .A2(n4659), .B1(N2873), .B2(n4693), .C1(n4742), 
        .C2(n7206), .Z(N4355) );
  AO222D0BWP U7977 ( .A1(N562), .A2(n4659), .B1(N2872), .B2(n4693), .C1(n4742), 
        .C2(n7207), .Z(N4354) );
  AO222D0BWP U7978 ( .A1(N561), .A2(n4659), .B1(N2871), .B2(n4693), .C1(n4741), 
        .C2(n7208), .Z(N4353) );
  AO222D0BWP U7979 ( .A1(N560), .A2(n4660), .B1(N2870), .B2(n4693), .C1(n4741), 
        .C2(n7209), .Z(N4352) );
  AO222D0BWP U7980 ( .A1(N559), .A2(n4660), .B1(N2869), .B2(n4694), .C1(n4741), 
        .C2(n7210), .Z(N4351) );
  AO222D0BWP U7981 ( .A1(N558), .A2(n4660), .B1(N2868), .B2(n4694), .C1(n4741), 
        .C2(n7211), .Z(N4350) );
  AO222D0BWP U7982 ( .A1(N557), .A2(n4660), .B1(N2867), .B2(n4694), .C1(n4741), 
        .C2(n7212), .Z(N4349) );
  AO222D0BWP U7983 ( .A1(N556), .A2(n4660), .B1(N2866), .B2(n4694), .C1(n4741), 
        .C2(n7213), .Z(N4348) );
  AO222D0BWP U7984 ( .A1(N555), .A2(n4660), .B1(N2865), .B2(n4694), .C1(n4741), 
        .C2(n7214), .Z(N4347) );
  AO222D0BWP U7985 ( .A1(N554), .A2(n4660), .B1(N2864), .B2(n4694), .C1(n4741), 
        .C2(n7215), .Z(N4346) );
  AO222D0BWP U7986 ( .A1(N553), .A2(n4660), .B1(N2863), .B2(n4694), .C1(n4741), 
        .C2(n7216), .Z(N4345) );
  AO222D0BWP U7987 ( .A1(N552), .A2(n4660), .B1(N2862), .B2(n4694), .C1(n4741), 
        .C2(n7217), .Z(N4344) );
  AO222D0BWP U7988 ( .A1(N551), .A2(n4660), .B1(N2861), .B2(n4694), .C1(n4741), 
        .C2(n7218), .Z(N4343) );
  AO222D0BWP U7989 ( .A1(N550), .A2(n4660), .B1(N2860), .B2(n4694), .C1(n4741), 
        .C2(n7219), .Z(N4342) );
  AO222D0BWP U7990 ( .A1(N549), .A2(n4660), .B1(N2859), .B2(n4694), .C1(n4740), 
        .C2(n7220), .Z(N4341) );
  AO222D0BWP U7991 ( .A1(N548), .A2(n4661), .B1(N2858), .B2(n4694), .C1(n4740), 
        .C2(n7221), .Z(N4340) );
  AO222D0BWP U7992 ( .A1(N547), .A2(n4661), .B1(N2857), .B2(n4694), .C1(n4740), 
        .C2(n7222), .Z(N4339) );
  AO222D0BWP U7993 ( .A1(N546), .A2(n4661), .B1(N2856), .B2(n4695), .C1(n4740), 
        .C2(n7223), .Z(N4338) );
  AO222D0BWP U7994 ( .A1(N545), .A2(n4661), .B1(N2855), .B2(n4695), .C1(n4740), 
        .C2(n7224), .Z(N4337) );
  AO222D0BWP U7995 ( .A1(N544), .A2(n4661), .B1(N2854), .B2(n4695), .C1(n4740), 
        .C2(n7225), .Z(N4336) );
  AO222D0BWP U7996 ( .A1(N543), .A2(n4661), .B1(N2853), .B2(n4695), .C1(n4740), 
        .C2(n7226), .Z(N4335) );
  AO222D0BWP U7997 ( .A1(N542), .A2(n4661), .B1(N2852), .B2(n4695), .C1(n4740), 
        .C2(n7227), .Z(N4334) );
  AO222D0BWP U7998 ( .A1(N541), .A2(n4661), .B1(N2851), .B2(n4695), .C1(n4740), 
        .C2(n7228), .Z(N4333) );
  AO222D0BWP U7999 ( .A1(N540), .A2(n4661), .B1(N2850), .B2(n4695), .C1(n4740), 
        .C2(n7229), .Z(N4332) );
  AO222D0BWP U8000 ( .A1(N539), .A2(n4661), .B1(N2849), .B2(n4695), .C1(n4740), 
        .C2(n7230), .Z(N4331) );
  AO222D0BWP U8001 ( .A1(N538), .A2(n4661), .B1(N2848), .B2(n4695), .C1(n4740), 
        .C2(n7231), .Z(N4330) );
  AO222D0BWP U8002 ( .A1(N537), .A2(n4661), .B1(N2847), .B2(n4695), .C1(n4739), 
        .C2(n7232), .Z(N4329) );
  AO222D0BWP U8003 ( .A1(N536), .A2(n4662), .B1(N2846), .B2(n4695), .C1(n4739), 
        .C2(n7233), .Z(N4328) );
  AO222D0BWP U8004 ( .A1(N535), .A2(n4662), .B1(N2845), .B2(n4695), .C1(n4739), 
        .C2(n7234), .Z(N4327) );
  AO222D0BWP U8005 ( .A1(N534), .A2(n4662), .B1(N2844), .B2(n4695), .C1(n4739), 
        .C2(n7235), .Z(N4326) );
  AO222D0BWP U8006 ( .A1(N533), .A2(n4662), .B1(N2843), .B2(n4696), .C1(n4739), 
        .C2(n7236), .Z(N4325) );
  AO222D0BWP U8007 ( .A1(N532), .A2(n4662), .B1(N2842), .B2(n4696), .C1(n4739), 
        .C2(n7237), .Z(N4324) );
  AO222D0BWP U8008 ( .A1(N531), .A2(n4662), .B1(N2841), .B2(n4696), .C1(n4739), 
        .C2(n7238), .Z(N4323) );
  OAI211D0BWP U8009 ( .A1(n6197), .A2(n6196), .B(n6204), .C(n6205), .ZN(N4322)
         );
  AO222D0BWP U8010 ( .A1(N530), .A2(n4662), .B1(N2840), .B2(n4696), .C1(n4739), 
        .C2(n7239), .Z(N4321) );
  AO222D0BWP U8011 ( .A1(N529), .A2(n4662), .B1(N2839), .B2(n4696), .C1(n4739), 
        .C2(n7240), .Z(N4320) );
  AO222D0BWP U8012 ( .A1(N528), .A2(n4662), .B1(N2838), .B2(n4696), .C1(n4739), 
        .C2(n7241), .Z(N4319) );
  AO222D0BWP U8013 ( .A1(N527), .A2(n4662), .B1(N2837), .B2(n4696), .C1(n4739), 
        .C2(n7242), .Z(N4318) );
  AO222D0BWP U8014 ( .A1(N526), .A2(n4662), .B1(N2836), .B2(n4696), .C1(n4739), 
        .C2(n7243), .Z(N4317) );
  AO222D0BWP U8015 ( .A1(N525), .A2(n4662), .B1(N2835), .B2(n4696), .C1(n4738), 
        .C2(n7244), .Z(N4316) );
  AO222D0BWP U8016 ( .A1(N524), .A2(n4663), .B1(N2834), .B2(n4696), .C1(n4738), 
        .C2(n7245), .Z(N4315) );
  AO222D0BWP U8017 ( .A1(N523), .A2(n4663), .B1(N2833), .B2(n4696), .C1(n4738), 
        .C2(n7246), .Z(N4314) );
  AO222D0BWP U8018 ( .A1(N522), .A2(n4663), .B1(N2832), .B2(n4696), .C1(n4738), 
        .C2(n7247), .Z(N4313) );
  AO222D0BWP U8019 ( .A1(N521), .A2(n4663), .B1(N2831), .B2(n4696), .C1(n4738), 
        .C2(n7248), .Z(N4312) );
  AO222D0BWP U8020 ( .A1(N520), .A2(n4663), .B1(N2830), .B2(n4697), .C1(n4738), 
        .C2(n7249), .Z(N4311) );
  AO222D0BWP U8021 ( .A1(N519), .A2(n4663), .B1(N2829), .B2(n4697), .C1(n4738), 
        .C2(n7250), .Z(N4310) );
  AO222D0BWP U8022 ( .A1(N518), .A2(n4663), .B1(N2828), .B2(n4697), .C1(n4738), 
        .C2(n7251), .Z(N4309) );
  AO222D0BWP U8023 ( .A1(N517), .A2(n4663), .B1(N2827), .B2(n4697), .C1(n4738), 
        .C2(n7252), .Z(N4308) );
  AO222D0BWP U8024 ( .A1(N516), .A2(n4663), .B1(N2826), .B2(n4697), .C1(n4738), 
        .C2(n7253), .Z(N4307) );
  AO222D0BWP U8025 ( .A1(N515), .A2(n4663), .B1(N2825), .B2(n4697), .C1(n4738), 
        .C2(n7254), .Z(N4306) );
  AO222D0BWP U8026 ( .A1(N514), .A2(n4663), .B1(N2824), .B2(n4697), .C1(n4738), 
        .C2(n7255), .Z(N4305) );
  AO222D0BWP U8027 ( .A1(N513), .A2(n4663), .B1(N2823), .B2(n4697), .C1(n4737), 
        .C2(n7256), .Z(N4304) );
  AO222D0BWP U8028 ( .A1(N512), .A2(n4664), .B1(N2822), .B2(n4697), .C1(n4737), 
        .C2(n7257), .Z(N4303) );
  AO222D0BWP U8029 ( .A1(N511), .A2(n4664), .B1(N2821), .B2(n4697), .C1(n4737), 
        .C2(n7258), .Z(N4302) );
  AO222D0BWP U8030 ( .A1(N510), .A2(n4664), .B1(N2820), .B2(n4697), .C1(n4737), 
        .C2(n7259), .Z(N4301) );
  AO222D0BWP U8031 ( .A1(N509), .A2(n4664), .B1(N2819), .B2(n4697), .C1(n4737), 
        .C2(n7260), .Z(N4300) );
  AO222D0BWP U8032 ( .A1(N508), .A2(n4664), .B1(N2818), .B2(n4697), .C1(n4737), 
        .C2(n7261), .Z(N4299) );
  AO222D0BWP U8033 ( .A1(N507), .A2(n4664), .B1(N2817), .B2(n4698), .C1(n4737), 
        .C2(n7262), .Z(N4298) );
  AO222D0BWP U8034 ( .A1(N506), .A2(n4664), .B1(N2816), .B2(n4698), .C1(n4737), 
        .C2(n7263), .Z(N4297) );
  AO222D0BWP U8035 ( .A1(N505), .A2(n4664), .B1(N2815), .B2(n4698), .C1(n4737), 
        .C2(n7264), .Z(N4296) );
  AO222D0BWP U8036 ( .A1(N504), .A2(n4664), .B1(N2814), .B2(n4698), .C1(n4737), 
        .C2(n7265), .Z(N4295) );
  AO222D0BWP U8037 ( .A1(N503), .A2(n4664), .B1(N2813), .B2(n4698), .C1(n4737), 
        .C2(n7266), .Z(N4294) );
  AO222D0BWP U8038 ( .A1(N502), .A2(n4664), .B1(N2812), .B2(n4698), .C1(n4737), 
        .C2(n7267), .Z(N4293) );
  AO222D0BWP U8039 ( .A1(N501), .A2(n4664), .B1(N2811), .B2(n4698), .C1(n4736), 
        .C2(n7268), .Z(N4292) );
  AO222D0BWP U8040 ( .A1(N500), .A2(n4665), .B1(N2810), .B2(n4698), .C1(n4736), 
        .C2(n7269), .Z(N4291) );
  AO222D0BWP U8041 ( .A1(N499), .A2(n4665), .B1(N2809), .B2(n4698), .C1(n4736), 
        .C2(n7270), .Z(N4290) );
  AO222D0BWP U8042 ( .A1(N498), .A2(n4665), .B1(N2808), .B2(n4698), .C1(n4736), 
        .C2(n7271), .Z(N4289) );
  AO222D0BWP U8043 ( .A1(N497), .A2(n4665), .B1(N2807), .B2(n4698), .C1(n4736), 
        .C2(n7272), .Z(N4288) );
  AO222D0BWP U8044 ( .A1(N496), .A2(n4665), .B1(N2806), .B2(n4698), .C1(n4736), 
        .C2(n7273), .Z(N4287) );
  AO222D0BWP U8045 ( .A1(N495), .A2(n4665), .B1(N2805), .B2(n4698), .C1(n4736), 
        .C2(n7274), .Z(N4286) );
  AO222D0BWP U8046 ( .A1(N494), .A2(n4665), .B1(N2804), .B2(n4699), .C1(n4736), 
        .C2(n7275), .Z(N4285) );
  AO222D0BWP U8047 ( .A1(N493), .A2(n4665), .B1(N2803), .B2(n4699), .C1(n4736), 
        .C2(n7276), .Z(N4284) );
  AO222D0BWP U8048 ( .A1(N492), .A2(n4665), .B1(N2802), .B2(n4699), .C1(n4736), 
        .C2(n7277), .Z(N4283) );
  AO222D0BWP U8049 ( .A1(N491), .A2(n4665), .B1(N2801), .B2(n4699), .C1(n4736), 
        .C2(n7278), .Z(N4282) );
  AO222D0BWP U8050 ( .A1(N490), .A2(n4665), .B1(N2800), .B2(n4699), .C1(n4736), 
        .C2(n7279), .Z(N4281) );
  AO222D0BWP U8051 ( .A1(N489), .A2(n4665), .B1(N2799), .B2(n4699), .C1(n4735), 
        .C2(n7280), .Z(N4280) );
  AO222D0BWP U8052 ( .A1(N488), .A2(n4666), .B1(N2798), .B2(n4699), .C1(n4735), 
        .C2(n7281), .Z(N4279) );
  AO222D0BWP U8053 ( .A1(N487), .A2(n4666), .B1(N2797), .B2(n4699), .C1(n4735), 
        .C2(n7282), .Z(N4278) );
  AO222D0BWP U8054 ( .A1(N486), .A2(n4666), .B1(N2796), .B2(n4699), .C1(n4735), 
        .C2(n7283), .Z(N4277) );
  AO222D0BWP U8055 ( .A1(N485), .A2(n4666), .B1(N2795), .B2(n4699), .C1(n4735), 
        .C2(n7284), .Z(N4276) );
  AO222D0BWP U8056 ( .A1(N484), .A2(n4666), .B1(N2794), .B2(n4699), .C1(n4735), 
        .C2(n7285), .Z(N4275) );
  AO222D0BWP U8057 ( .A1(N483), .A2(n4666), .B1(N2793), .B2(n4699), .C1(n4735), 
        .C2(n7286), .Z(N4274) );
  AO222D0BWP U8058 ( .A1(N482), .A2(n4666), .B1(N2792), .B2(n4699), .C1(n4735), 
        .C2(n7287), .Z(N4273) );
  AO222D0BWP U8059 ( .A1(N481), .A2(n4666), .B1(N2791), .B2(n4700), .C1(n4735), 
        .C2(n7288), .Z(N4272) );
  AO222D0BWP U8060 ( .A1(N480), .A2(n4666), .B1(N2790), .B2(n4700), .C1(n4735), 
        .C2(n7289), .Z(N4271) );
  AO222D0BWP U8061 ( .A1(N479), .A2(n4666), .B1(N2789), .B2(n4700), .C1(n4735), 
        .C2(n7290), .Z(N4270) );
  AO222D0BWP U8062 ( .A1(N478), .A2(n4666), .B1(N2788), .B2(n4700), .C1(n4735), 
        .C2(n7291), .Z(N4269) );
  AO222D0BWP U8063 ( .A1(N477), .A2(n4666), .B1(N2787), .B2(n4700), .C1(n4734), 
        .C2(n7292), .Z(N4268) );
  AO222D0BWP U8064 ( .A1(N476), .A2(n4667), .B1(N2786), .B2(n4700), .C1(n4734), 
        .C2(n7293), .Z(N4267) );
  AO222D0BWP U8065 ( .A1(N475), .A2(n4667), .B1(N2785), .B2(n4700), .C1(n4734), 
        .C2(n7294), .Z(N4266) );
  AO222D0BWP U8066 ( .A1(N474), .A2(n4667), .B1(N2784), .B2(n4700), .C1(n4734), 
        .C2(n7295), .Z(N4265) );
  AO222D0BWP U8067 ( .A1(N473), .A2(n4667), .B1(N2783), .B2(n4700), .C1(n4734), 
        .C2(n7296), .Z(N4264) );
  AO222D0BWP U8068 ( .A1(N472), .A2(n4667), .B1(N2782), .B2(n4700), .C1(n4734), 
        .C2(n7297), .Z(N4263) );
  AO222D0BWP U8069 ( .A1(N471), .A2(n4667), .B1(N2781), .B2(n4700), .C1(n4734), 
        .C2(n7298), .Z(N4262) );
  AO222D0BWP U8070 ( .A1(N470), .A2(n4667), .B1(N2780), .B2(n4700), .C1(n4734), 
        .C2(n7299), .Z(N4261) );
  AO222D0BWP U8071 ( .A1(N469), .A2(n4667), .B1(N2779), .B2(n4700), .C1(n4734), 
        .C2(n7300), .Z(N4260) );
  AO222D0BWP U8072 ( .A1(N468), .A2(n4667), .B1(N2778), .B2(n4701), .C1(n4734), 
        .C2(n7301), .Z(N4259) );
  AO222D0BWP U8073 ( .A1(N467), .A2(n4667), .B1(N2777), .B2(n4701), .C1(n4734), 
        .C2(n7302), .Z(N4258) );
  AO222D0BWP U8074 ( .A1(N466), .A2(n4667), .B1(N2776), .B2(n4701), .C1(n4734), 
        .C2(n7303), .Z(N4257) );
  AO222D0BWP U8075 ( .A1(N465), .A2(n4667), .B1(N2775), .B2(n4701), .C1(n4733), 
        .C2(n7304), .Z(N4256) );
  AO222D0BWP U8076 ( .A1(N464), .A2(n4668), .B1(N2774), .B2(n4701), .C1(n4733), 
        .C2(n7305), .Z(N4255) );
  AO222D0BWP U8077 ( .A1(N463), .A2(n4668), .B1(N2773), .B2(n4701), .C1(n4733), 
        .C2(n7306), .Z(N4254) );
  AO222D0BWP U8078 ( .A1(N462), .A2(n4668), .B1(N2772), .B2(n4701), .C1(n4733), 
        .C2(n7307), .Z(N4253) );
  AO222D0BWP U8079 ( .A1(N461), .A2(n4668), .B1(N2771), .B2(n4701), .C1(n4733), 
        .C2(n7308), .Z(N4252) );
  AO222D0BWP U8080 ( .A1(N460), .A2(n4668), .B1(N2770), .B2(n4701), .C1(n4733), 
        .C2(n7309), .Z(N4251) );
  AO222D0BWP U8081 ( .A1(N459), .A2(n4668), .B1(N2769), .B2(n4701), .C1(n4733), 
        .C2(n7310), .Z(N4250) );
  AO222D0BWP U8082 ( .A1(N458), .A2(n4668), .B1(N2768), .B2(n4701), .C1(n4733), 
        .C2(n7311), .Z(N4249) );
  AO222D0BWP U8083 ( .A1(N457), .A2(n4668), .B1(N2767), .B2(n4701), .C1(n4733), 
        .C2(n7312), .Z(N4248) );
  AO222D0BWP U8084 ( .A1(N456), .A2(n4668), .B1(N2766), .B2(n4701), .C1(n4733), 
        .C2(n7313), .Z(N4247) );
  AO222D0BWP U8085 ( .A1(N455), .A2(n4668), .B1(N2765), .B2(n4702), .C1(n4733), 
        .C2(n7314), .Z(N4246) );
  AO222D0BWP U8086 ( .A1(N454), .A2(n4668), .B1(N2764), .B2(n4702), .C1(n4733), 
        .C2(n7315), .Z(N4245) );
  AO222D0BWP U8087 ( .A1(N453), .A2(n4668), .B1(N2763), .B2(n4702), .C1(n4732), 
        .C2(n7316), .Z(N4244) );
  AO222D0BWP U8088 ( .A1(N452), .A2(n4669), .B1(N2762), .B2(n4702), .C1(n4732), 
        .C2(n7317), .Z(N4243) );
  AO222D0BWP U8089 ( .A1(N451), .A2(n4669), .B1(N2761), .B2(n4702), .C1(n4732), 
        .C2(n7318), .Z(N4242) );
  AO222D0BWP U8090 ( .A1(N450), .A2(n4669), .B1(N2760), .B2(n4702), .C1(n4732), 
        .C2(n7319), .Z(N4241) );
  AO222D0BWP U8091 ( .A1(N449), .A2(n4669), .B1(N2759), .B2(n4702), .C1(n4732), 
        .C2(n7320), .Z(N4240) );
  AO222D0BWP U8092 ( .A1(N448), .A2(n4669), .B1(N2758), .B2(n4702), .C1(n4732), 
        .C2(n7321), .Z(N4239) );
  AO222D0BWP U8093 ( .A1(N447), .A2(n4669), .B1(N2757), .B2(n4702), .C1(n4732), 
        .C2(n7322), .Z(N4238) );
  AO222D0BWP U8094 ( .A1(N446), .A2(n4669), .B1(N2756), .B2(n4702), .C1(n4732), 
        .C2(n7323), .Z(N4237) );
  AO222D0BWP U8095 ( .A1(N445), .A2(n4669), .B1(N2755), .B2(n4702), .C1(n4732), 
        .C2(n7324), .Z(N4236) );
  AO222D0BWP U8096 ( .A1(N444), .A2(n4669), .B1(N2754), .B2(n4702), .C1(n4732), 
        .C2(n7325), .Z(N4235) );
  AO222D0BWP U8097 ( .A1(N443), .A2(n4669), .B1(N2753), .B2(n4702), .C1(n4732), 
        .C2(n7326), .Z(N4234) );
  AO222D0BWP U8098 ( .A1(N442), .A2(n4669), .B1(N2752), .B2(n4703), .C1(n4732), 
        .C2(n7327), .Z(N4233) );
  AO222D0BWP U8099 ( .A1(N441), .A2(n4669), .B1(N2751), .B2(n4703), .C1(n4731), 
        .C2(n7328), .Z(N4232) );
  AO222D0BWP U8100 ( .A1(N440), .A2(n4670), .B1(N2750), .B2(n4703), .C1(n4731), 
        .C2(n7329), .Z(N4231) );
  AO222D0BWP U8101 ( .A1(N439), .A2(n4670), .B1(N2749), .B2(n4703), .C1(n4731), 
        .C2(n7330), .Z(N4230) );
  AO222D0BWP U8102 ( .A1(N438), .A2(n4670), .B1(N2748), .B2(n4703), .C1(n4731), 
        .C2(n7331), .Z(N4229) );
  AO222D0BWP U8103 ( .A1(N437), .A2(n4670), .B1(N2747), .B2(n4703), .C1(n4731), 
        .C2(n7332), .Z(N4228) );
  AO222D0BWP U8104 ( .A1(N436), .A2(n4670), .B1(N2746), .B2(n4703), .C1(n4731), 
        .C2(n7333), .Z(N4227) );
  AO222D0BWP U8105 ( .A1(N435), .A2(n4670), .B1(N2745), .B2(n4703), .C1(n4731), 
        .C2(n7334), .Z(N4226) );
  AO222D0BWP U8106 ( .A1(N434), .A2(n4670), .B1(N2744), .B2(n4703), .C1(n4731), 
        .C2(n7335), .Z(N4225) );
  AO222D0BWP U8107 ( .A1(N433), .A2(n4670), .B1(N2743), .B2(n4703), .C1(n4731), 
        .C2(n7336), .Z(N4224) );
  AO222D0BWP U8108 ( .A1(N432), .A2(n4670), .B1(N2742), .B2(n4703), .C1(n4731), 
        .C2(n7337), .Z(N4223) );
  AO222D0BWP U8109 ( .A1(N431), .A2(n4670), .B1(N2741), .B2(n4703), .C1(n4731), 
        .C2(n7338), .Z(N4221) );
  AO222D0BWP U8110 ( .A1(N430), .A2(n4670), .B1(N2740), .B2(n4703), .C1(n4731), 
        .C2(n7339), .Z(N4220) );
  AO222D0BWP U8111 ( .A1(N429), .A2(n4670), .B1(N2739), .B2(n4704), .C1(n4730), 
        .C2(n7340), .Z(N4219) );
  AO222D0BWP U8112 ( .A1(N428), .A2(n4671), .B1(N2738), .B2(n4704), .C1(n4730), 
        .C2(n7341), .Z(N4218) );
  AO222D0BWP U8113 ( .A1(N427), .A2(n4671), .B1(N2737), .B2(n4704), .C1(n4730), 
        .C2(n7342), .Z(N4217) );
  AO222D0BWP U8114 ( .A1(N426), .A2(n4671), .B1(N2736), .B2(n4704), .C1(n4730), 
        .C2(n7343), .Z(N4216) );
  AO222D0BWP U8115 ( .A1(N425), .A2(n4671), .B1(N2735), .B2(n4704), .C1(n4730), 
        .C2(n7344), .Z(N4215) );
  AO222D0BWP U8116 ( .A1(N424), .A2(n4671), .B1(N2734), .B2(n4704), .C1(n4730), 
        .C2(n7345), .Z(N4214) );
  AO222D0BWP U8117 ( .A1(N423), .A2(n4671), .B1(N2733), .B2(n4704), .C1(n4730), 
        .C2(n7346), .Z(N4213) );
  AO222D0BWP U8118 ( .A1(N422), .A2(n4671), .B1(N2732), .B2(n4704), .C1(n4730), 
        .C2(n7347), .Z(N4212) );
  AO222D0BWP U8119 ( .A1(N421), .A2(n4671), .B1(N2731), .B2(n4704), .C1(n4730), 
        .C2(n7348), .Z(N4211) );
  AO222D0BWP U8120 ( .A1(N420), .A2(n4671), .B1(N2730), .B2(n4704), .C1(n4730), 
        .C2(n7349), .Z(N4210) );
  AO222D0BWP U8121 ( .A1(N419), .A2(n4671), .B1(N2729), .B2(n4704), .C1(n4730), 
        .C2(n7350), .Z(N4209) );
  AO222D0BWP U8122 ( .A1(N418), .A2(n4671), .B1(N2728), .B2(n4704), .C1(n4730), 
        .C2(n7351), .Z(N4208) );
  AO222D0BWP U8123 ( .A1(N417), .A2(n4671), .B1(N2727), .B2(n4704), .C1(n4729), 
        .C2(n7352), .Z(N4207) );
  AO222D0BWP U8124 ( .A1(N416), .A2(n4672), .B1(N2726), .B2(n4705), .C1(n4729), 
        .C2(n7353), .Z(N4206) );
  AO222D0BWP U8125 ( .A1(N415), .A2(n4672), .B1(N2725), .B2(n4705), .C1(n4729), 
        .C2(n7354), .Z(N4205) );
  AO222D0BWP U8126 ( .A1(N414), .A2(n4672), .B1(N2724), .B2(n4705), .C1(n4729), 
        .C2(n7355), .Z(N4204) );
  AO222D0BWP U8127 ( .A1(N413), .A2(n4672), .B1(N2723), .B2(n4705), .C1(n4729), 
        .C2(n7356), .Z(N4203) );
  AO222D0BWP U8128 ( .A1(N412), .A2(n4672), .B1(N2722), .B2(n4705), .C1(n4729), 
        .C2(n7357), .Z(N4202) );
  AO222D0BWP U8129 ( .A1(N411), .A2(n4672), .B1(N2721), .B2(n4705), .C1(n4729), 
        .C2(n7358), .Z(N4201) );
  AO222D0BWP U8130 ( .A1(N410), .A2(n4672), .B1(N2720), .B2(n4705), .C1(n4729), 
        .C2(n7359), .Z(N4200) );
  AO222D0BWP U8131 ( .A1(N409), .A2(n4672), .B1(N2719), .B2(n4705), .C1(n4729), 
        .C2(n7360), .Z(N4199) );
  AO222D0BWP U8132 ( .A1(N408), .A2(n4672), .B1(N2718), .B2(n4705), .C1(n4729), 
        .C2(n7361), .Z(N4198) );
  AO222D0BWP U8133 ( .A1(N407), .A2(n4672), .B1(N2717), .B2(n4705), .C1(n4729), 
        .C2(n7362), .Z(N4197) );
  AO222D0BWP U8134 ( .A1(N406), .A2(n4672), .B1(N2716), .B2(n4705), .C1(n4729), 
        .C2(n7363), .Z(N4196) );
  AO222D0BWP U8135 ( .A1(N405), .A2(n4672), .B1(N2715), .B2(n4705), .C1(n4728), 
        .C2(n7364), .Z(N4195) );
  AO222D0BWP U8136 ( .A1(N404), .A2(n4673), .B1(N2714), .B2(n4705), .C1(n4728), 
        .C2(n7365), .Z(N4194) );
  AO222D0BWP U8137 ( .A1(N403), .A2(n4673), .B1(N2713), .B2(n4706), .C1(n4728), 
        .C2(n7366), .Z(N4193) );
  AO222D0BWP U8138 ( .A1(N402), .A2(n4673), .B1(N2712), .B2(n4706), .C1(n4728), 
        .C2(n7367), .Z(N4192) );
  AO222D0BWP U8139 ( .A1(N401), .A2(n4673), .B1(N2711), .B2(n4706), .C1(n4728), 
        .C2(n7368), .Z(N4191) );
  AO222D0BWP U8140 ( .A1(N400), .A2(n4673), .B1(N2710), .B2(n4706), .C1(n4728), 
        .C2(n7369), .Z(N4190) );
  AO222D0BWP U8141 ( .A1(N399), .A2(n4673), .B1(N2709), .B2(n4706), .C1(n4728), 
        .C2(n7370), .Z(N4189) );
  AO222D0BWP U8142 ( .A1(N398), .A2(n4673), .B1(N2708), .B2(n4706), .C1(n4728), 
        .C2(n7371), .Z(N4188) );
  AO222D0BWP U8143 ( .A1(N397), .A2(n4673), .B1(N2707), .B2(n4706), .C1(n4728), 
        .C2(n7372), .Z(N4187) );
  AO222D0BWP U8144 ( .A1(N396), .A2(n4673), .B1(N2706), .B2(n4706), .C1(n4728), 
        .C2(n7373), .Z(N4186) );
  AO222D0BWP U8145 ( .A1(N395), .A2(n4673), .B1(N2705), .B2(n4706), .C1(n4728), 
        .C2(n7374), .Z(N4185) );
  AO222D0BWP U8146 ( .A1(N394), .A2(n4673), .B1(N2704), .B2(n4706), .C1(n4728), 
        .C2(n7375), .Z(N4184) );
  AO222D0BWP U8147 ( .A1(N393), .A2(n4673), .B1(N2703), .B2(n4706), .C1(n4727), 
        .C2(n7376), .Z(N4183) );
  AO222D0BWP U8148 ( .A1(N392), .A2(n4674), .B1(N2702), .B2(n4706), .C1(n4727), 
        .C2(n7377), .Z(N4182) );
  AO222D0BWP U8149 ( .A1(N391), .A2(n4674), .B1(N2701), .B2(n4706), .C1(n4727), 
        .C2(n7378), .Z(N4181) );
  AO222D0BWP U8150 ( .A1(N390), .A2(n4674), .B1(N2700), .B2(n4707), .C1(n4727), 
        .C2(n7379), .Z(N4180) );
  AO222D0BWP U8151 ( .A1(N389), .A2(n4674), .B1(N2699), .B2(n4707), .C1(n4727), 
        .C2(n7380), .Z(N4179) );
  AO222D0BWP U8152 ( .A1(N388), .A2(n4674), .B1(N2698), .B2(n4707), .C1(n4727), 
        .C2(n7381), .Z(N4178) );
  AO222D0BWP U8153 ( .A1(N387), .A2(n4674), .B1(N2697), .B2(n4707), .C1(n4727), 
        .C2(n7382), .Z(N4177) );
  AO222D0BWP U8154 ( .A1(N386), .A2(n4674), .B1(N2696), .B2(n4707), .C1(n4727), 
        .C2(n7383), .Z(N4176) );
  AO222D0BWP U8155 ( .A1(N385), .A2(n4674), .B1(N2695), .B2(n4707), .C1(n4727), 
        .C2(n7384), .Z(N4175) );
  AO222D0BWP U8156 ( .A1(N384), .A2(n4674), .B1(N2694), .B2(n4707), .C1(n4727), 
        .C2(n7385), .Z(N4174) );
  AO222D0BWP U8157 ( .A1(N383), .A2(n4674), .B1(N2693), .B2(n4707), .C1(n4727), 
        .C2(n7386), .Z(N4173) );
  AO222D0BWP U8158 ( .A1(N382), .A2(n4674), .B1(N2692), .B2(n4707), .C1(n4727), 
        .C2(n7387), .Z(N4172) );
  AO222D0BWP U8159 ( .A1(N381), .A2(n4674), .B1(N2691), .B2(n4707), .C1(n4726), 
        .C2(n7388), .Z(N4171) );
  AO222D0BWP U8160 ( .A1(N380), .A2(n4675), .B1(N2690), .B2(n4707), .C1(n4726), 
        .C2(n7389), .Z(N4170) );
  AO222D0BWP U8161 ( .A1(N379), .A2(n4675), .B1(N2689), .B2(n4707), .C1(n4726), 
        .C2(n7390), .Z(N4169) );
  AO222D0BWP U8162 ( .A1(N378), .A2(n4675), .B1(N2688), .B2(n4707), .C1(n4726), 
        .C2(n7391), .Z(N4168) );
  AO222D0BWP U8163 ( .A1(N377), .A2(n4675), .B1(N2687), .B2(n4708), .C1(n4726), 
        .C2(n7392), .Z(N4167) );
  AO222D0BWP U8164 ( .A1(N376), .A2(n4675), .B1(N2686), .B2(n4708), .C1(n4726), 
        .C2(n7393), .Z(N4166) );
  AO222D0BWP U8165 ( .A1(N375), .A2(n4675), .B1(N2685), .B2(n4708), .C1(n4726), 
        .C2(n7394), .Z(N4165) );
  AO222D0BWP U8166 ( .A1(N374), .A2(n4675), .B1(N2684), .B2(n4708), .C1(n4726), 
        .C2(n7395), .Z(N4164) );
  AO222D0BWP U8167 ( .A1(N373), .A2(n4675), .B1(N2683), .B2(n4708), .C1(n4726), 
        .C2(n7396), .Z(N4163) );
  AO222D0BWP U8168 ( .A1(N372), .A2(n4675), .B1(N2682), .B2(n4708), .C1(n4726), 
        .C2(n7397), .Z(N4162) );
  AO222D0BWP U8169 ( .A1(N371), .A2(n4675), .B1(N2681), .B2(n4708), .C1(n4726), 
        .C2(n7398), .Z(N4161) );
  AO222D0BWP U8170 ( .A1(N370), .A2(n4675), .B1(N2680), .B2(n4708), .C1(n4726), 
        .C2(n7399), .Z(N4160) );
  AO222D0BWP U8171 ( .A1(N369), .A2(n4675), .B1(N2679), .B2(n4708), .C1(n4725), 
        .C2(n7400), .Z(N4159) );
  AO222D0BWP U8172 ( .A1(N368), .A2(n4676), .B1(N2678), .B2(n4708), .C1(n4725), 
        .C2(n7401), .Z(N4158) );
  AO222D0BWP U8173 ( .A1(N367), .A2(n4676), .B1(N2677), .B2(n4708), .C1(n4725), 
        .C2(n7402), .Z(N4157) );
  AO222D0BWP U8174 ( .A1(N366), .A2(n4676), .B1(N2676), .B2(n4708), .C1(n4725), 
        .C2(n7403), .Z(N4156) );
  AO222D0BWP U8175 ( .A1(N365), .A2(n4676), .B1(N2675), .B2(n4708), .C1(n4725), 
        .C2(n7404), .Z(N4155) );
  AO222D0BWP U8176 ( .A1(N364), .A2(n4676), .B1(N2674), .B2(n4709), .C1(n4725), 
        .C2(n7405), .Z(N4154) );
  AO222D0BWP U8177 ( .A1(N363), .A2(n4676), .B1(N2673), .B2(n4709), .C1(n4725), 
        .C2(n7406), .Z(N4153) );
  AO222D0BWP U8178 ( .A1(N362), .A2(n4676), .B1(N2672), .B2(n4709), .C1(n4725), 
        .C2(n7407), .Z(N4152) );
  AO222D0BWP U8179 ( .A1(N361), .A2(n4676), .B1(N2671), .B2(n4709), .C1(n4725), 
        .C2(n7408), .Z(N4151) );
  AO222D0BWP U8180 ( .A1(N360), .A2(n4676), .B1(N2670), .B2(n4709), .C1(n4725), 
        .C2(n7409), .Z(N4150) );
  AO222D0BWP U8181 ( .A1(N359), .A2(n4676), .B1(N2669), .B2(n4709), .C1(n4725), 
        .C2(n7410), .Z(N4149) );
  AO222D0BWP U8182 ( .A1(N358), .A2(n4676), .B1(N2668), .B2(n4709), .C1(n4725), 
        .C2(n7411), .Z(N4148) );
  AO222D0BWP U8183 ( .A1(N357), .A2(n4676), .B1(N2667), .B2(n4709), .C1(n4724), 
        .C2(n7412), .Z(N4147) );
  AO222D0BWP U8184 ( .A1(N356), .A2(n4677), .B1(N2666), .B2(n4709), .C1(n4724), 
        .C2(n7413), .Z(N4146) );
  AO222D0BWP U8185 ( .A1(N355), .A2(n4677), .B1(N2665), .B2(n4709), .C1(n4724), 
        .C2(n7414), .Z(N4145) );
  AO222D0BWP U8186 ( .A1(N354), .A2(n4677), .B1(N2664), .B2(n4709), .C1(n4724), 
        .C2(n7415), .Z(N4144) );
  AO222D0BWP U8187 ( .A1(N353), .A2(n4677), .B1(N2663), .B2(n4709), .C1(n4724), 
        .C2(n7416), .Z(N4143) );
  AO222D0BWP U8188 ( .A1(N352), .A2(n4677), .B1(N2662), .B2(n4709), .C1(n4724), 
        .C2(n7417), .Z(N4142) );
  AO222D0BWP U8189 ( .A1(N351), .A2(n4677), .B1(N2661), .B2(n4710), .C1(n4724), 
        .C2(n7418), .Z(N4141) );
  AO222D0BWP U8190 ( .A1(N350), .A2(n4677), .B1(N2660), .B2(n4710), .C1(n4724), 
        .C2(n7419), .Z(N4140) );
  AO222D0BWP U8191 ( .A1(N349), .A2(n4677), .B1(N2659), .B2(n4710), .C1(n4724), 
        .C2(n7420), .Z(N4139) );
  AO222D0BWP U8192 ( .A1(N348), .A2(n4677), .B1(N2658), .B2(n4710), .C1(n4724), 
        .C2(n7421), .Z(N4138) );
  AO222D0BWP U8193 ( .A1(N347), .A2(n4677), .B1(N2657), .B2(n4710), .C1(n4724), 
        .C2(n7422), .Z(N4137) );
  AO222D0BWP U8194 ( .A1(N346), .A2(n4677), .B1(N2656), .B2(n4710), .C1(n4724), 
        .C2(n7423), .Z(N4136) );
  AO222D0BWP U8195 ( .A1(N345), .A2(n4677), .B1(N2655), .B2(n4710), .C1(n4723), 
        .C2(n7424), .Z(N4135) );
  AO222D0BWP U8196 ( .A1(N344), .A2(n4678), .B1(N2654), .B2(n4710), .C1(n4723), 
        .C2(n7425), .Z(N4134) );
  AO222D0BWP U8197 ( .A1(N343), .A2(n4678), .B1(N2653), .B2(n4710), .C1(n4723), 
        .C2(n7426), .Z(N4133) );
  AO222D0BWP U8198 ( .A1(N342), .A2(n4678), .B1(N2652), .B2(n4710), .C1(n4723), 
        .C2(n7427), .Z(N4132) );
  AO222D0BWP U8199 ( .A1(N341), .A2(n4678), .B1(N2651), .B2(n4710), .C1(n4723), 
        .C2(n7428), .Z(N4131) );
  AO222D0BWP U8200 ( .A1(N340), .A2(n4678), .B1(N2650), .B2(n4710), .C1(n4723), 
        .C2(n7429), .Z(N4130) );
  AO222D0BWP U8201 ( .A1(N339), .A2(n4678), .B1(N2649), .B2(n4710), .C1(n4723), 
        .C2(n7430), .Z(N4129) );
  AO222D0BWP U8202 ( .A1(N338), .A2(n4678), .B1(N2648), .B2(n4711), .C1(n4723), 
        .C2(n7431), .Z(N4128) );
  AO222D0BWP U8203 ( .A1(N337), .A2(n4678), .B1(N2647), .B2(n4711), .C1(n4723), 
        .C2(n7432), .Z(N4127) );
  AO222D0BWP U8204 ( .A1(N336), .A2(n4678), .B1(N2646), .B2(n4711), .C1(n4723), 
        .C2(n7433), .Z(N4126) );
  AO222D0BWP U8205 ( .A1(N335), .A2(n4678), .B1(N2645), .B2(n4711), .C1(n4723), 
        .C2(n7434), .Z(N4125) );
  AO222D0BWP U8206 ( .A1(N334), .A2(n4678), .B1(N2644), .B2(n4711), .C1(n4723), 
        .C2(n7435), .Z(N4124) );
  CKND0BWP U8207 ( .I(n6206), .ZN(n6203) );
  OAI211D0BWP U8208 ( .A1(n3419), .A2(n6206), .B(n6207), .C(n6208), .ZN(N4123)
         );
  AOI32D0BWP U8209 ( .A1(n6209), .A2(n6210), .A3(n7476), .B1(N2643), .B2(n4711), .ZN(n6208) );
  CKND0BWP U8210 ( .I(n6211), .ZN(n7476) );
  CKND2D0BWP U8211 ( .A1(N333), .A2(n4678), .ZN(n6207) );
  OAI211D0BWP U8212 ( .A1(n3403), .A2(n6206), .B(n6212), .C(n6213), .ZN(N4121)
         );
  AOI222D0BWP U8213 ( .A1(DataIn[15]), .A2(n6214), .B1(N2642), .B2(n6215), 
        .C1(n6216), .C2(result[15]), .ZN(n6213) );
  CKND2D0BWP U8214 ( .A1(N332), .A2(n4678), .ZN(n6212) );
  OAI211D0BWP U8215 ( .A1(n3404), .A2(n6206), .B(n6217), .C(n6218), .ZN(N4120)
         );
  AOI222D0BWP U8216 ( .A1(DataIn[14]), .A2(n6214), .B1(N2641), .B2(n6215), 
        .C1(n6216), .C2(result[14]), .ZN(n6218) );
  CKND2D0BWP U8217 ( .A1(N331), .A2(n4679), .ZN(n6217) );
  OAI211D0BWP U8218 ( .A1(n3405), .A2(n6206), .B(n6219), .C(n6220), .ZN(N4119)
         );
  AOI222D0BWP U8219 ( .A1(DataIn[13]), .A2(n6214), .B1(N2640), .B2(n6215), 
        .C1(n6216), .C2(result[13]), .ZN(n6220) );
  CKND2D0BWP U8220 ( .A1(N330), .A2(n4679), .ZN(n6219) );
  OAI211D0BWP U8221 ( .A1(n3406), .A2(n6206), .B(n6221), .C(n6222), .ZN(N4118)
         );
  AOI222D0BWP U8222 ( .A1(DataIn[12]), .A2(n6214), .B1(N2639), .B2(n6215), 
        .C1(n6216), .C2(result[12]), .ZN(n6222) );
  CKND2D0BWP U8223 ( .A1(N329), .A2(n4679), .ZN(n6221) );
  OAI211D0BWP U8224 ( .A1(n3407), .A2(n6206), .B(n6223), .C(n6224), .ZN(N4117)
         );
  AOI222D0BWP U8225 ( .A1(DataIn[11]), .A2(n6214), .B1(N2638), .B2(n6215), 
        .C1(n6216), .C2(result[11]), .ZN(n6224) );
  CKND2D0BWP U8226 ( .A1(N328), .A2(n4679), .ZN(n6223) );
  OAI211D0BWP U8227 ( .A1(n3408), .A2(n6206), .B(n6225), .C(n6226), .ZN(N4116)
         );
  AOI222D0BWP U8228 ( .A1(DataIn[10]), .A2(n6214), .B1(N2637), .B2(n6215), 
        .C1(n6216), .C2(result[10]), .ZN(n6226) );
  CKND2D0BWP U8229 ( .A1(N327), .A2(n4679), .ZN(n6225) );
  OAI211D0BWP U8230 ( .A1(n3409), .A2(n6206), .B(n6227), .C(n6228), .ZN(N4115)
         );
  AOI222D0BWP U8231 ( .A1(DataIn[9]), .A2(n6214), .B1(N2636), .B2(n6215), .C1(
        n6216), .C2(result[9]), .ZN(n6228) );
  CKND2D0BWP U8232 ( .A1(N326), .A2(n4679), .ZN(n6227) );
  OAI211D0BWP U8233 ( .A1(n3410), .A2(n6206), .B(n6229), .C(n6230), .ZN(N4114)
         );
  AOI222D0BWP U8234 ( .A1(DataIn[8]), .A2(n6214), .B1(N2635), .B2(n6215), .C1(
        n6216), .C2(result[8]), .ZN(n6230) );
  CKND2D0BWP U8235 ( .A1(N325), .A2(n4679), .ZN(n6229) );
  OAI211D0BWP U8236 ( .A1(n3411), .A2(n6206), .B(n6231), .C(n6232), .ZN(N4113)
         );
  AOI222D0BWP U8237 ( .A1(DataIn[7]), .A2(n6214), .B1(N2634), .B2(n6215), .C1(
        n6216), .C2(result[7]), .ZN(n6232) );
  CKND2D0BWP U8238 ( .A1(N324), .A2(n4679), .ZN(n6231) );
  OAI211D0BWP U8239 ( .A1(n3412), .A2(n6206), .B(n6233), .C(n6234), .ZN(N4112)
         );
  AOI222D0BWP U8240 ( .A1(DataIn[6]), .A2(n6214), .B1(N2633), .B2(n6215), .C1(
        n6216), .C2(result[6]), .ZN(n6234) );
  CKND2D0BWP U8241 ( .A1(N323), .A2(n4679), .ZN(n6233) );
  OAI211D0BWP U8242 ( .A1(n3413), .A2(n6206), .B(n6235), .C(n6236), .ZN(N4111)
         );
  AOI222D0BWP U8243 ( .A1(DataIn[5]), .A2(n6214), .B1(N2632), .B2(n6215), .C1(
        n6216), .C2(result[5]), .ZN(n6236) );
  CKND2D0BWP U8244 ( .A1(N322), .A2(n4679), .ZN(n6235) );
  OAI211D0BWP U8245 ( .A1(n3414), .A2(n6206), .B(n6237), .C(n6238), .ZN(N4110)
         );
  AOI222D0BWP U8246 ( .A1(DataIn[4]), .A2(n6214), .B1(N2631), .B2(n6215), .C1(
        n6216), .C2(result[4]), .ZN(n6238) );
  CKND2D0BWP U8247 ( .A1(N321), .A2(n4679), .ZN(n6237) );
  OAI211D0BWP U8248 ( .A1(n3415), .A2(n6206), .B(n6239), .C(n6240), .ZN(N4109)
         );
  AOI222D0BWP U8249 ( .A1(DataIn[3]), .A2(n6214), .B1(N2630), .B2(n6215), .C1(
        n6216), .C2(result[3]), .ZN(n6240) );
  CKND2D0BWP U8250 ( .A1(N320), .A2(n4679), .ZN(n6239) );
  OAI211D0BWP U8251 ( .A1(n3416), .A2(n6206), .B(n6241), .C(n6242), .ZN(N4108)
         );
  AOI222D0BWP U8252 ( .A1(DataIn[2]), .A2(n6214), .B1(N2629), .B2(n6215), .C1(
        n6216), .C2(result[2]), .ZN(n6242) );
  CKND2D0BWP U8253 ( .A1(N319), .A2(n4679), .ZN(n6241) );
  OAI211D0BWP U8254 ( .A1(n3417), .A2(n6206), .B(n6243), .C(n6244), .ZN(N4107)
         );
  AOI222D0BWP U8255 ( .A1(DataIn[1]), .A2(n6214), .B1(N2628), .B2(n6215), .C1(
        n6216), .C2(result[1]), .ZN(n6244) );
  CKND2D0BWP U8256 ( .A1(N318), .A2(n4680), .ZN(n6243) );
  OAI211D0BWP U8257 ( .A1(n3418), .A2(n6206), .B(n6245), .C(n6246), .ZN(N4106)
         );
  AOI222D0BWP U8258 ( .A1(DataIn[0]), .A2(n6214), .B1(N2627), .B2(n6215), .C1(
        n6216), .C2(result[0]), .ZN(n6246) );
  NR2D0BWP U8259 ( .A1(n6196), .A2(n6205), .ZN(n6216) );
  INR2D0BWP U8260 ( .A1(n4711), .B1(n5988), .ZN(n6214) );
  NR2D0BWP U8261 ( .A1(n6197), .A2(n6210), .ZN(n6202) );
  CKND2D0BWP U8262 ( .A1(N317), .A2(n4680), .ZN(n6245) );
  NR2D0BWP U8263 ( .A1(n6210), .A2(n6205), .ZN(n6201) );
  CKND2D0BWP U8264 ( .A1(N4105), .A2(n6196), .ZN(n6206) );
  OAI31D0BWP U8265 ( .A1(n6247), .A2(n6248), .A3(n6249), .B(n6250), .ZN(N4103)
         );
  ND3D0BWP U8266 ( .A1(N4104), .A2(n6211), .A3(n6251), .ZN(n6249) );
  OAI211D0BWP U8267 ( .A1(op1[15]), .A2(n5963), .B(n6252), .C(n6253), .ZN(
        n6211) );
  NR2D0BWP U8268 ( .A1(n6254), .A2(n6255), .ZN(n6253) );
  MUX2ND0BWP U8269 ( .I0(n5485), .I1(n6256), .S(n6121), .ZN(n6255) );
  NR2D0BWP U8270 ( .A1(func[2]), .A2(func[1]), .ZN(n6121) );
  MUX2ND0BWP U8271 ( .I0(n6257), .I1(n6122), .S(func[2]), .ZN(n6254) );
  CKND0BWP U8272 ( .I(func[1]), .ZN(n6122) );
  CKND2D0BWP U8273 ( .A1(n6256), .A2(n5485), .ZN(n6257) );
  CKND0BWP U8274 ( .I(func[0]), .ZN(n6256) );
  AO21D0BWP U8275 ( .A1(n5963), .A2(op1[15]), .B(op2[15]), .Z(n6252) );
  OAI22D0BWP U8276 ( .A1(n5964), .A2(n5965), .B1(n6258), .B2(n6005), .ZN(n5963) );
  CKND0BWP U8277 ( .I(op2[14]), .ZN(n6005) );
  NR2D0BWP U8278 ( .A1(\alu/N851 ), .A2(n6259), .ZN(n6258) );
  CKND0BWP U8279 ( .I(\alu/N851 ), .ZN(n5965) );
  CKND0BWP U8280 ( .I(n6259), .ZN(n5964) );
  OAI22D0BWP U8281 ( .A1(n5966), .A2(n5967), .B1(n6260), .B2(n6030), .ZN(n6259) );
  CKND0BWP U8282 ( .I(op2[13]), .ZN(n6030) );
  NR2D0BWP U8283 ( .A1(op1[13]), .A2(n6261), .ZN(n6260) );
  CKND0BWP U8284 ( .I(op1[13]), .ZN(n5967) );
  CKND0BWP U8285 ( .I(n6261), .ZN(n5966) );
  OAI22D0BWP U8286 ( .A1(n5968), .A2(n5969), .B1(n6262), .B2(n6036), .ZN(n6261) );
  CKND0BWP U8287 ( .I(op2[12]), .ZN(n6036) );
  NR2D0BWP U8288 ( .A1(op1[12]), .A2(n6263), .ZN(n6262) );
  CKND0BWP U8289 ( .I(op1[12]), .ZN(n5969) );
  CKND0BWP U8290 ( .I(n6263), .ZN(n5968) );
  OAI22D0BWP U8291 ( .A1(n5970), .A2(n5971), .B1(n6264), .B2(n6015), .ZN(n6263) );
  CKND0BWP U8292 ( .I(op2[11]), .ZN(n6015) );
  NR2D0BWP U8293 ( .A1(op1[11]), .A2(n6265), .ZN(n6264) );
  CKND0BWP U8294 ( .I(op1[11]), .ZN(n5971) );
  CKND0BWP U8295 ( .I(n6265), .ZN(n5970) );
  OAI22D0BWP U8296 ( .A1(n5972), .A2(n5973), .B1(n6266), .B2(n6018), .ZN(n6265) );
  CKND0BWP U8297 ( .I(op2[10]), .ZN(n6018) );
  NR2D0BWP U8298 ( .A1(op1[10]), .A2(n6267), .ZN(n6266) );
  CKND0BWP U8299 ( .I(op1[10]), .ZN(n5973) );
  CKND0BWP U8300 ( .I(n6267), .ZN(n5972) );
  OAI22D0BWP U8301 ( .A1(n5974), .A2(n5975), .B1(n6268), .B2(n6045), .ZN(n6267) );
  CKND0BWP U8302 ( .I(op2[9]), .ZN(n6045) );
  NR2D0BWP U8303 ( .A1(op1[9]), .A2(n6269), .ZN(n6268) );
  CKND0BWP U8304 ( .I(op1[9]), .ZN(n5975) );
  CKND0BWP U8305 ( .I(n6269), .ZN(n5974) );
  OAI22D0BWP U8306 ( .A1(n5976), .A2(n5977), .B1(n6270), .B2(n6046), .ZN(n6269) );
  CKND0BWP U8307 ( .I(op2[8]), .ZN(n6046) );
  NR2D0BWP U8308 ( .A1(op1[8]), .A2(n6271), .ZN(n6270) );
  CKND0BWP U8309 ( .I(op1[8]), .ZN(n5977) );
  CKND0BWP U8310 ( .I(n6271), .ZN(n5976) );
  OAI22D0BWP U8311 ( .A1(n5978), .A2(n3370), .B1(n6272), .B2(n3374), .ZN(n6271) );
  AN2D0BWP U8312 ( .A1(n5978), .A2(n3370), .Z(n6272) );
  MAOI22D0BWP U8313 ( .A1(n5979), .A2(op1[6]), .B1(n6273), .B2(n3372), .ZN(
        n5978) );
  NR2D0BWP U8314 ( .A1(op1[6]), .A2(n5979), .ZN(n6273) );
  MOAI22D0BWP U8315 ( .A1(n6274), .A2(n3378), .B1(n5980), .B2(op1[5]), .ZN(
        n5979) );
  NR2D0BWP U8316 ( .A1(op1[5]), .A2(n5980), .ZN(n6274) );
  MOAI22D0BWP U8317 ( .A1(n6275), .A2(n3373), .B1(n5981), .B2(op1[4]), .ZN(
        n5980) );
  NR2D0BWP U8318 ( .A1(op1[4]), .A2(n5981), .ZN(n6275) );
  MOAI22D0BWP U8319 ( .A1(n6276), .A2(n3375), .B1(n5982), .B2(op1[3]), .ZN(
        n5981) );
  NR2D0BWP U8320 ( .A1(op1[3]), .A2(n5982), .ZN(n6276) );
  OAI22D0BWP U8321 ( .A1(n6277), .A2(n3371), .B1(n6278), .B2(n3379), .ZN(n5982) );
  NR2D0BWP U8322 ( .A1(op1[2]), .A2(n5983), .ZN(n6278) );
  CKND0BWP U8323 ( .I(n6277), .ZN(n5983) );
  MAOI222D0BWP U8324 ( .A(op2[1]), .B(op1[1]), .C(n6279), .ZN(n6277) );
  NR2D0BWP U8325 ( .A1(n6048), .A2(n6047), .ZN(n6279) );
  CKND0BWP U8326 ( .I(op2[0]), .ZN(n6047) );
  CKND0BWP U8327 ( .I(op1[0]), .ZN(n6048) );
  ND4D0BWP U8328 ( .A1(n5998), .A2(n6186), .A3(n5997), .A4(n5996), .ZN(n6248)
         );
  ND4D0BWP U8329 ( .A1(n5994), .A2(n5993), .A3(n5995), .A4(n6280), .ZN(n6247)
         );
  NR4D0BWP U8330 ( .A1(result[9]), .A2(result[8]), .A3(result[7]), .A4(
        result[6]), .ZN(n6280) );
  CKND2D0BWP U8331 ( .A1(n6205), .A2(n2522), .ZN(N4104) );
  OAI211D0BWP U8332 ( .A1(n3645), .A2(n6281), .B(n6282), .C(n6283), .ZN(N4101)
         );
  AOI22D0BWP U8333 ( .A1(n6199), .A2(n6284), .B1(n6285), .B2(scalarData2[15]), 
        .ZN(n6283) );
  ND4D0BWP U8334 ( .A1(n6286), .A2(n6287), .A3(n6288), .A4(n6289), .ZN(n6284)
         );
  AOI221D0BWP U8335 ( .A1(vectorData2[159]), .A2(n6290), .B1(vectorData2[175]), 
        .B2(n6291), .C(n6292), .ZN(n6289) );
  MOAI22D0BWP U8336 ( .A1(n6293), .A2(n3546), .B1(n6294), .B2(vectorData2[143]), .ZN(n6292) );
  AOI221D0BWP U8337 ( .A1(vectorData2[207]), .A2(n6295), .B1(vectorData2[223]), 
        .B2(n6296), .C(n6297), .ZN(n6288) );
  OAI22D0BWP U8338 ( .A1(n6298), .A2(n3498), .B1(n6299), .B2(n3600), .ZN(n6297) );
  AOI221D0BWP U8339 ( .A1(vectorData2[47]), .A2(n6300), .B1(vectorData2[63]), 
        .B2(n6301), .C(n6302), .ZN(n6287) );
  AO22D0BWP U8340 ( .A1(n6303), .A2(vectorData2[255]), .B1(n6304), .B2(
        vectorData2[239]), .Z(n6302) );
  AOI222D0BWP U8341 ( .A1(vectorData2[111]), .A2(n6305), .B1(vectorData2[79]), 
        .B2(n6306), .C1(vectorData2[95]), .C2(n6307), .ZN(n6286) );
  OAI211D0BWP U8342 ( .A1(n3642), .A2(n6281), .B(n6282), .C(n6308), .ZN(N4100)
         );
  AOI22D0BWP U8343 ( .A1(n6199), .A2(n6309), .B1(n6285), .B2(scalarData2[14]), 
        .ZN(n6308) );
  ND4D0BWP U8344 ( .A1(n6310), .A2(n6311), .A3(n6312), .A4(n6313), .ZN(n6309)
         );
  AOI221D0BWP U8345 ( .A1(vectorData2[158]), .A2(n6290), .B1(vectorData2[174]), 
        .B2(n6291), .C(n6314), .ZN(n6313) );
  MOAI22D0BWP U8346 ( .A1(n6293), .A2(n3543), .B1(n6294), .B2(vectorData2[142]), .ZN(n6314) );
  AOI221D0BWP U8347 ( .A1(vectorData2[206]), .A2(n6295), .B1(vectorData2[222]), 
        .B2(n6296), .C(n6315), .ZN(n6312) );
  OAI22D0BWP U8348 ( .A1(n6298), .A2(n3495), .B1(n6299), .B2(n3597), .ZN(n6315) );
  AOI221D0BWP U8349 ( .A1(vectorData2[46]), .A2(n6300), .B1(vectorData2[62]), 
        .B2(n6301), .C(n6316), .ZN(n6311) );
  AO22D0BWP U8350 ( .A1(n6303), .A2(vectorData2[254]), .B1(n6304), .B2(
        vectorData2[238]), .Z(n6316) );
  AOI222D0BWP U8351 ( .A1(vectorData2[110]), .A2(n6305), .B1(vectorData2[78]), 
        .B2(n6306), .C1(vectorData2[94]), .C2(n6307), .ZN(n6310) );
  OAI211D0BWP U8352 ( .A1(n3639), .A2(n6281), .B(n6282), .C(n6317), .ZN(N4099)
         );
  AOI22D0BWP U8353 ( .A1(n6199), .A2(n6318), .B1(n6285), .B2(scalarData2[13]), 
        .ZN(n6317) );
  ND4D0BWP U8354 ( .A1(n6319), .A2(n6320), .A3(n6321), .A4(n6322), .ZN(n6318)
         );
  AOI221D0BWP U8355 ( .A1(vectorData2[157]), .A2(n6290), .B1(vectorData2[173]), 
        .B2(n6291), .C(n6323), .ZN(n6322) );
  MOAI22D0BWP U8356 ( .A1(n6293), .A2(n3540), .B1(n6294), .B2(vectorData2[141]), .ZN(n6323) );
  AOI221D0BWP U8357 ( .A1(vectorData2[205]), .A2(n6295), .B1(vectorData2[221]), 
        .B2(n6296), .C(n6324), .ZN(n6321) );
  OAI22D0BWP U8358 ( .A1(n6298), .A2(n3492), .B1(n6299), .B2(n3594), .ZN(n6324) );
  AOI221D0BWP U8359 ( .A1(vectorData2[45]), .A2(n6300), .B1(vectorData2[61]), 
        .B2(n6301), .C(n6325), .ZN(n6320) );
  AO22D0BWP U8360 ( .A1(n6303), .A2(vectorData2[253]), .B1(n6304), .B2(
        vectorData2[237]), .Z(n6325) );
  AOI222D0BWP U8361 ( .A1(vectorData2[109]), .A2(n6305), .B1(vectorData2[77]), 
        .B2(n6306), .C1(vectorData2[93]), .C2(n6307), .ZN(n6319) );
  OAI211D0BWP U8362 ( .A1(n3636), .A2(n6281), .B(n6282), .C(n6326), .ZN(N4098)
         );
  AOI22D0BWP U8363 ( .A1(n6199), .A2(n6327), .B1(n6285), .B2(scalarData2[12]), 
        .ZN(n6326) );
  ND4D0BWP U8364 ( .A1(n6328), .A2(n6329), .A3(n6330), .A4(n6331), .ZN(n6327)
         );
  AOI221D0BWP U8365 ( .A1(vectorData2[156]), .A2(n6290), .B1(vectorData2[172]), 
        .B2(n6291), .C(n6332), .ZN(n6331) );
  MOAI22D0BWP U8366 ( .A1(n6293), .A2(n3537), .B1(n6294), .B2(vectorData2[140]), .ZN(n6332) );
  AOI221D0BWP U8367 ( .A1(vectorData2[204]), .A2(n6295), .B1(vectorData2[220]), 
        .B2(n6296), .C(n6333), .ZN(n6330) );
  OAI22D0BWP U8368 ( .A1(n6298), .A2(n3489), .B1(n6299), .B2(n3591), .ZN(n6333) );
  AOI221D0BWP U8369 ( .A1(vectorData2[44]), .A2(n6300), .B1(vectorData2[60]), 
        .B2(n6301), .C(n6334), .ZN(n6329) );
  AO22D0BWP U8370 ( .A1(n6303), .A2(vectorData2[252]), .B1(n6304), .B2(
        vectorData2[236]), .Z(n6334) );
  AOI222D0BWP U8371 ( .A1(vectorData2[108]), .A2(n6305), .B1(vectorData2[76]), 
        .B2(n6306), .C1(vectorData2[92]), .C2(n6307), .ZN(n6328) );
  OAI211D0BWP U8372 ( .A1(n3633), .A2(n6281), .B(n6282), .C(n6335), .ZN(N4097)
         );
  AOI22D0BWP U8373 ( .A1(n6199), .A2(n6336), .B1(n6285), .B2(scalarData2[11]), 
        .ZN(n6335) );
  ND4D0BWP U8374 ( .A1(n6337), .A2(n6338), .A3(n6339), .A4(n6340), .ZN(n6336)
         );
  AOI221D0BWP U8375 ( .A1(vectorData2[155]), .A2(n6290), .B1(vectorData2[171]), 
        .B2(n6291), .C(n6341), .ZN(n6340) );
  MOAI22D0BWP U8376 ( .A1(n6293), .A2(n3534), .B1(n6294), .B2(vectorData2[139]), .ZN(n6341) );
  AOI221D0BWP U8377 ( .A1(vectorData2[203]), .A2(n6295), .B1(vectorData2[219]), 
        .B2(n6296), .C(n6342), .ZN(n6339) );
  OAI22D0BWP U8378 ( .A1(n6298), .A2(n3486), .B1(n6299), .B2(n3588), .ZN(n6342) );
  AOI221D0BWP U8379 ( .A1(vectorData2[43]), .A2(n6300), .B1(vectorData2[59]), 
        .B2(n6301), .C(n6343), .ZN(n6338) );
  AO22D0BWP U8380 ( .A1(n6303), .A2(vectorData2[251]), .B1(n6304), .B2(
        vectorData2[235]), .Z(n6343) );
  AOI222D0BWP U8381 ( .A1(vectorData2[107]), .A2(n6305), .B1(vectorData2[75]), 
        .B2(n6306), .C1(vectorData2[91]), .C2(n6307), .ZN(n6337) );
  AOI21D0BWP U8382 ( .A1(instrIn[11]), .A2(n6344), .B(n6345), .ZN(n6282) );
  OAI221D0BWP U8383 ( .A1(n3699), .A2(n6346), .B1(n3672), .B2(n6281), .C(n6347), .ZN(N4096) );
  AOI221D0BWP U8384 ( .A1(n6199), .A2(n6348), .B1(n6344), .B2(instrIn[10]), 
        .C(n6345), .ZN(n6347) );
  ND4D0BWP U8385 ( .A1(n6349), .A2(n6350), .A3(n6351), .A4(n6352), .ZN(n6348)
         );
  AOI221D0BWP U8386 ( .A1(vectorData2[154]), .A2(n6290), .B1(vectorData2[170]), 
        .B2(n6291), .C(n6353), .ZN(n6352) );
  MOAI22D0BWP U8387 ( .A1(n6293), .A2(n3531), .B1(n6294), .B2(vectorData2[138]), .ZN(n6353) );
  AOI221D0BWP U8388 ( .A1(vectorData2[202]), .A2(n6295), .B1(vectorData2[218]), 
        .B2(n6296), .C(n6354), .ZN(n6351) );
  OAI22D0BWP U8389 ( .A1(n6298), .A2(n3483), .B1(n6299), .B2(n3585), .ZN(n6354) );
  AOI221D0BWP U8390 ( .A1(vectorData2[42]), .A2(n6300), .B1(vectorData2[58]), 
        .B2(n6301), .C(n6355), .ZN(n6350) );
  AO22D0BWP U8391 ( .A1(n6303), .A2(vectorData2[250]), .B1(n6304), .B2(
        vectorData2[234]), .Z(n6355) );
  AOI222D0BWP U8392 ( .A1(vectorData2[106]), .A2(n6305), .B1(vectorData2[74]), 
        .B2(n6306), .C1(vectorData2[90]), .C2(n6307), .ZN(n6349) );
  OAI221D0BWP U8393 ( .A1(n3696), .A2(n6346), .B1(n3669), .B2(n6281), .C(n6356), .ZN(N4095) );
  AOI221D0BWP U8394 ( .A1(n6199), .A2(n6357), .B1(n6344), .B2(instrIn[9]), .C(
        n6345), .ZN(n6356) );
  ND4D0BWP U8395 ( .A1(n6358), .A2(n6359), .A3(n6360), .A4(n6361), .ZN(n6357)
         );
  AOI221D0BWP U8396 ( .A1(vectorData2[153]), .A2(n6290), .B1(vectorData2[169]), 
        .B2(n6291), .C(n6362), .ZN(n6361) );
  MOAI22D0BWP U8397 ( .A1(n6293), .A2(n3528), .B1(n6294), .B2(vectorData2[137]), .ZN(n6362) );
  AOI221D0BWP U8398 ( .A1(vectorData2[201]), .A2(n6295), .B1(vectorData2[217]), 
        .B2(n6296), .C(n6363), .ZN(n6360) );
  OAI22D0BWP U8399 ( .A1(n6298), .A2(n3480), .B1(n6299), .B2(n3582), .ZN(n6363) );
  AOI221D0BWP U8400 ( .A1(vectorData2[41]), .A2(n6300), .B1(vectorData2[57]), 
        .B2(n6301), .C(n6364), .ZN(n6359) );
  AO22D0BWP U8401 ( .A1(n6303), .A2(vectorData2[249]), .B1(n6304), .B2(
        vectorData2[233]), .Z(n6364) );
  AOI222D0BWP U8402 ( .A1(vectorData2[105]), .A2(n6305), .B1(vectorData2[73]), 
        .B2(n6306), .C1(vectorData2[89]), .C2(n6307), .ZN(n6358) );
  OAI221D0BWP U8403 ( .A1(n3693), .A2(n6346), .B1(n3666), .B2(n6281), .C(n6365), .ZN(N4094) );
  AOI221D0BWP U8404 ( .A1(n6199), .A2(n6366), .B1(n6344), .B2(instrIn[8]), .C(
        n6345), .ZN(n6365) );
  ND4D0BWP U8405 ( .A1(n6367), .A2(n6368), .A3(n6369), .A4(n6370), .ZN(n6366)
         );
  AOI221D0BWP U8406 ( .A1(vectorData2[152]), .A2(n6290), .B1(vectorData2[168]), 
        .B2(n6291), .C(n6371), .ZN(n6370) );
  MOAI22D0BWP U8407 ( .A1(n6293), .A2(n3525), .B1(n6294), .B2(vectorData2[136]), .ZN(n6371) );
  AOI221D0BWP U8408 ( .A1(vectorData2[200]), .A2(n6295), .B1(vectorData2[216]), 
        .B2(n6296), .C(n6372), .ZN(n6369) );
  OAI22D0BWP U8409 ( .A1(n6298), .A2(n3477), .B1(n6299), .B2(n3579), .ZN(n6372) );
  AOI221D0BWP U8410 ( .A1(vectorData2[40]), .A2(n6300), .B1(vectorData2[56]), 
        .B2(n6301), .C(n6373), .ZN(n6368) );
  AO22D0BWP U8411 ( .A1(n6303), .A2(vectorData2[248]), .B1(n6304), .B2(
        vectorData2[232]), .Z(n6373) );
  AOI222D0BWP U8412 ( .A1(vectorData2[104]), .A2(n6305), .B1(vectorData2[72]), 
        .B2(n6306), .C1(vectorData2[88]), .C2(n6307), .ZN(n6367) );
  OAI221D0BWP U8413 ( .A1(n3690), .A2(n6346), .B1(n3663), .B2(n6281), .C(n6374), .ZN(N4093) );
  AOI221D0BWP U8414 ( .A1(instrIn[7]), .A2(n6375), .B1(n6199), .B2(n6376), .C(
        n6345), .ZN(n6374) );
  ND4D0BWP U8415 ( .A1(n6377), .A2(n6378), .A3(n6379), .A4(n6380), .ZN(n6376)
         );
  AOI221D0BWP U8416 ( .A1(vectorData2[151]), .A2(n6290), .B1(vectorData2[167]), 
        .B2(n6291), .C(n6381), .ZN(n6380) );
  MOAI22D0BWP U8417 ( .A1(n6293), .A2(n3558), .B1(n6294), .B2(vectorData2[135]), .ZN(n6381) );
  AOI221D0BWP U8418 ( .A1(vectorData2[199]), .A2(n6295), .B1(vectorData2[215]), 
        .B2(n6296), .C(n6382), .ZN(n6379) );
  OAI22D0BWP U8419 ( .A1(n6298), .A2(n3510), .B1(n6299), .B2(n3612), .ZN(n6382) );
  AOI221D0BWP U8420 ( .A1(vectorData2[39]), .A2(n6300), .B1(vectorData2[55]), 
        .B2(n6301), .C(n6383), .ZN(n6378) );
  AO22D0BWP U8421 ( .A1(n6303), .A2(vectorData2[247]), .B1(n6304), .B2(
        vectorData2[231]), .Z(n6383) );
  AOI222D0BWP U8422 ( .A1(vectorData2[103]), .A2(n6305), .B1(vectorData2[71]), 
        .B2(n6306), .C1(vectorData2[87]), .C2(n6307), .ZN(n6377) );
  OAI221D0BWP U8423 ( .A1(n3687), .A2(n6346), .B1(n3660), .B2(n6281), .C(n6384), .ZN(N4092) );
  AOI221D0BWP U8424 ( .A1(instrIn[6]), .A2(n6375), .B1(n6199), .B2(n6385), .C(
        n6345), .ZN(n6384) );
  ND4D0BWP U8425 ( .A1(n6386), .A2(n6387), .A3(n6388), .A4(n6389), .ZN(n6385)
         );
  AOI221D0BWP U8426 ( .A1(vectorData2[150]), .A2(n6290), .B1(vectorData2[166]), 
        .B2(n6291), .C(n6390), .ZN(n6389) );
  MOAI22D0BWP U8427 ( .A1(n6293), .A2(n3555), .B1(n6294), .B2(vectorData2[134]), .ZN(n6390) );
  AOI221D0BWP U8428 ( .A1(vectorData2[198]), .A2(n6295), .B1(vectorData2[214]), 
        .B2(n6296), .C(n6391), .ZN(n6388) );
  OAI22D0BWP U8429 ( .A1(n6298), .A2(n3507), .B1(n6299), .B2(n3609), .ZN(n6391) );
  AOI221D0BWP U8430 ( .A1(vectorData2[38]), .A2(n6300), .B1(vectorData2[54]), 
        .B2(n6301), .C(n6392), .ZN(n6387) );
  AO22D0BWP U8431 ( .A1(n6303), .A2(vectorData2[246]), .B1(n6304), .B2(
        vectorData2[230]), .Z(n6392) );
  AOI222D0BWP U8432 ( .A1(vectorData2[102]), .A2(n6305), .B1(vectorData2[70]), 
        .B2(n6306), .C1(vectorData2[86]), .C2(n6307), .ZN(n6386) );
  OAI221D0BWP U8433 ( .A1(n3684), .A2(n6346), .B1(n3657), .B2(n6281), .C(n6393), .ZN(N4091) );
  AOI221D0BWP U8434 ( .A1(instrIn[5]), .A2(n6375), .B1(n6199), .B2(n6394), .C(
        n6345), .ZN(n6393) );
  NR3D0BWP U8435 ( .A1(n6395), .A2(n6396), .A3(n5537), .ZN(n6345) );
  CKND0BWP U8436 ( .I(instrIn[5]), .ZN(n5537) );
  ND4D0BWP U8437 ( .A1(n6397), .A2(n6398), .A3(n6399), .A4(n6400), .ZN(n6394)
         );
  AOI221D0BWP U8438 ( .A1(vectorData2[149]), .A2(n6290), .B1(vectorData2[165]), 
        .B2(n6291), .C(n6401), .ZN(n6400) );
  MOAI22D0BWP U8439 ( .A1(n6293), .A2(n3552), .B1(n6294), .B2(vectorData2[133]), .ZN(n6401) );
  AOI221D0BWP U8440 ( .A1(vectorData2[197]), .A2(n6295), .B1(vectorData2[213]), 
        .B2(n6296), .C(n6402), .ZN(n6399) );
  OAI22D0BWP U8441 ( .A1(n6298), .A2(n3504), .B1(n6299), .B2(n3606), .ZN(n6402) );
  AOI221D0BWP U8442 ( .A1(vectorData2[37]), .A2(n6300), .B1(vectorData2[53]), 
        .B2(n6301), .C(n6403), .ZN(n6398) );
  AO22D0BWP U8443 ( .A1(n6303), .A2(vectorData2[245]), .B1(n6304), .B2(
        vectorData2[229]), .Z(n6403) );
  AOI222D0BWP U8444 ( .A1(vectorData2[101]), .A2(n6305), .B1(vectorData2[69]), 
        .B2(n6306), .C1(vectorData2[85]), .C2(n6307), .ZN(n6397) );
  CKND0BWP U8445 ( .I(n6404), .ZN(n6375) );
  OAI221D0BWP U8446 ( .A1(n6405), .A2(n6406), .B1(n6407), .B2(n5540), .C(n6408), .ZN(N4090) );
  AOI22D0BWP U8447 ( .A1(n6285), .A2(scalarData2[4]), .B1(n6409), .B2(
        vectorData2[4]), .ZN(n6408) );
  CKND0BWP U8448 ( .I(instrIn[4]), .ZN(n5540) );
  NR4D0BWP U8449 ( .A1(n6410), .A2(n6411), .A3(n6412), .A4(n6413), .ZN(n6405)
         );
  OAI222D0BWP U8450 ( .A1(n6414), .A2(n3516), .B1(n6415), .B2(n3624), .C1(
        n6416), .C2(n3618), .ZN(n6413) );
  OAI221D0BWP U8451 ( .A1(n6417), .A2(n3462), .B1(n6418), .B2(n3570), .C(n6419), .ZN(n6412) );
  AOI22D0BWP U8452 ( .A1(vectorData2[228]), .A2(n6304), .B1(vectorData2[244]), 
        .B2(n6303), .ZN(n6419) );
  OAI221D0BWP U8453 ( .A1(n6420), .A2(n3468), .B1(n6421), .B2(n3564), .C(n6422), .ZN(n6411) );
  AOI22D0BWP U8454 ( .A1(vectorData2[20]), .A2(n6423), .B1(vectorData2[180]), 
        .B2(n6424), .ZN(n6422) );
  OAI221D0BWP U8455 ( .A1(n6425), .A2(n6426), .B1(n6427), .B2(n3630), .C(n6428), .ZN(n6410) );
  AOI22D0BWP U8456 ( .A1(vectorData2[116]), .A2(n6429), .B1(vectorData2[132]), 
        .B2(n6294), .ZN(n6428) );
  CKND0BWP U8457 ( .I(vectorData2[148]), .ZN(n6426) );
  OAI221D0BWP U8458 ( .A1(n6430), .A2(n6406), .B1(n6407), .B2(n5542), .C(n6431), .ZN(N4089) );
  AOI22D0BWP U8459 ( .A1(n6285), .A2(scalarData2[3]), .B1(n6409), .B2(
        vectorData2[3]), .ZN(n6431) );
  CKND0BWP U8460 ( .I(instrIn[3]), .ZN(n5542) );
  CKND0BWP U8461 ( .I(n6432), .ZN(n6407) );
  NR4D0BWP U8462 ( .A1(n6433), .A2(n6434), .A3(n6435), .A4(n6436), .ZN(n6430)
         );
  OAI222D0BWP U8463 ( .A1(n6414), .A2(n3513), .B1(n6415), .B2(n3621), .C1(
        n6416), .C2(n3615), .ZN(n6436) );
  OAI221D0BWP U8464 ( .A1(n6417), .A2(n3459), .B1(n6418), .B2(n3567), .C(n6437), .ZN(n6435) );
  AOI22D0BWP U8465 ( .A1(vectorData2[227]), .A2(n6304), .B1(vectorData2[243]), 
        .B2(n6303), .ZN(n6437) );
  OAI221D0BWP U8466 ( .A1(n6420), .A2(n3465), .B1(n6421), .B2(n3561), .C(n6438), .ZN(n6434) );
  AOI22D0BWP U8467 ( .A1(vectorData2[19]), .A2(n6423), .B1(vectorData2[179]), 
        .B2(n6424), .ZN(n6438) );
  CKND0BWP U8468 ( .I(n6298), .ZN(n6424) );
  CKND0BWP U8469 ( .I(n6299), .ZN(n6423) );
  OAI221D0BWP U8470 ( .A1(n6425), .A2(n6439), .B1(n6427), .B2(n3627), .C(n6440), .ZN(n6433) );
  AOI22D0BWP U8471 ( .A1(vectorData2[115]), .A2(n6429), .B1(vectorData2[131]), 
        .B2(n6294), .ZN(n6440) );
  CKND0BWP U8472 ( .I(n6293), .ZN(n6429) );
  CKND0BWP U8473 ( .I(vectorData2[147]), .ZN(n6439) );
  OAI221D0BWP U8474 ( .A1(n3681), .A2(n6346), .B1(n3654), .B2(n6281), .C(n6441), .ZN(N4088) );
  AOI22D0BWP U8475 ( .A1(n6199), .A2(n6442), .B1(instrIn[2]), .B2(n6432), .ZN(
        n6441) );
  ND4D0BWP U8476 ( .A1(n6443), .A2(n6444), .A3(n6445), .A4(n6446), .ZN(n6442)
         );
  AOI221D0BWP U8477 ( .A1(vectorData2[146]), .A2(n6290), .B1(vectorData2[162]), 
        .B2(n6291), .C(n6447), .ZN(n6446) );
  MOAI22D0BWP U8478 ( .A1(n6293), .A2(n3549), .B1(n6294), .B2(vectorData2[130]), .ZN(n6447) );
  AOI221D0BWP U8479 ( .A1(vectorData2[194]), .A2(n6295), .B1(vectorData2[210]), 
        .B2(n6296), .C(n6448), .ZN(n6445) );
  OAI22D0BWP U8480 ( .A1(n6298), .A2(n3501), .B1(n6299), .B2(n3603), .ZN(n6448) );
  AOI221D0BWP U8481 ( .A1(vectorData2[34]), .A2(n6300), .B1(vectorData2[50]), 
        .B2(n6301), .C(n6449), .ZN(n6444) );
  AO22D0BWP U8482 ( .A1(n6303), .A2(vectorData2[242]), .B1(n6304), .B2(
        vectorData2[226]), .Z(n6449) );
  AOI222D0BWP U8483 ( .A1(vectorData2[98]), .A2(n6305), .B1(vectorData2[66]), 
        .B2(n6306), .C1(vectorData2[82]), .C2(n6307), .ZN(n6443) );
  OAI221D0BWP U8484 ( .A1(n3678), .A2(n6346), .B1(n3651), .B2(n6281), .C(n6450), .ZN(N4087) );
  AOI22D0BWP U8485 ( .A1(n6199), .A2(n6451), .B1(instrIn[1]), .B2(n6432), .ZN(
        n6450) );
  ND4D0BWP U8486 ( .A1(n6452), .A2(n6453), .A3(n6454), .A4(n6455), .ZN(n6451)
         );
  AOI221D0BWP U8487 ( .A1(vectorData2[145]), .A2(n6290), .B1(vectorData2[161]), 
        .B2(n6291), .C(n6456), .ZN(n6455) );
  MOAI22D0BWP U8488 ( .A1(n6293), .A2(n3522), .B1(n6294), .B2(vectorData2[129]), .ZN(n6456) );
  AOI221D0BWP U8489 ( .A1(vectorData2[193]), .A2(n6295), .B1(vectorData2[209]), 
        .B2(n6296), .C(n6457), .ZN(n6454) );
  OAI22D0BWP U8490 ( .A1(n6298), .A2(n3474), .B1(n6299), .B2(n3576), .ZN(n6457) );
  AOI221D0BWP U8491 ( .A1(vectorData2[33]), .A2(n6300), .B1(vectorData2[49]), 
        .B2(n6301), .C(n6458), .ZN(n6453) );
  AO22D0BWP U8492 ( .A1(n6303), .A2(vectorData2[241]), .B1(n6304), .B2(
        vectorData2[225]), .Z(n6458) );
  AOI222D0BWP U8493 ( .A1(vectorData2[97]), .A2(n6305), .B1(vectorData2[65]), 
        .B2(n6306), .C1(vectorData2[81]), .C2(n6307), .ZN(n6452) );
  OAI221D0BWP U8494 ( .A1(n3675), .A2(n6346), .B1(n3648), .B2(n6281), .C(n6459), .ZN(N4086) );
  AOI22D0BWP U8495 ( .A1(instrIn[0]), .A2(n6432), .B1(n6199), .B2(n6460), .ZN(
        n6459) );
  ND4D0BWP U8496 ( .A1(n6461), .A2(n6462), .A3(n6463), .A4(n6464), .ZN(n6460)
         );
  AOI221D0BWP U8497 ( .A1(vectorData2[144]), .A2(n6290), .B1(vectorData2[160]), 
        .B2(n6291), .C(n6465), .ZN(n6464) );
  MOAI22D0BWP U8498 ( .A1(n6293), .A2(n3519), .B1(n6294), .B2(vectorData2[128]), .ZN(n6465) );
  AO22D0BWP U8499 ( .A1(n6466), .A2(N1101), .B1(n6467), .B2(N260), .Z(n6294)
         );
  AOI22D0BWP U8500 ( .A1(n6466), .A2(N1100), .B1(n6467), .B2(N259), .ZN(n6293)
         );
  CKND0BWP U8501 ( .I(n6427), .ZN(n6291) );
  AOI22D0BWP U8502 ( .A1(n6466), .A2(N1103), .B1(n6467), .B2(N262), .ZN(n6427)
         );
  CKND0BWP U8503 ( .I(n6425), .ZN(n6290) );
  AOI22D0BWP U8504 ( .A1(n6466), .A2(N1102), .B1(n6467), .B2(N261), .ZN(n6425)
         );
  AOI221D0BWP U8505 ( .A1(vectorData2[192]), .A2(n6295), .B1(vectorData2[208]), 
        .B2(n6296), .C(n6468), .ZN(n6463) );
  OAI22D0BWP U8506 ( .A1(n6298), .A2(n3471), .B1(n6299), .B2(n3573), .ZN(n6468) );
  AOI22D0BWP U8507 ( .A1(n6466), .A2(N1094), .B1(n6467), .B2(N253), .ZN(n6299)
         );
  AOI22D0BWP U8508 ( .A1(n6466), .A2(N1104), .B1(n6467), .B2(N263), .ZN(n6298)
         );
  CKND0BWP U8509 ( .I(n6421), .ZN(n6296) );
  AOI22D0BWP U8510 ( .A1(n6466), .A2(N1106), .B1(n6467), .B2(N265), .ZN(n6421)
         );
  CKND0BWP U8511 ( .I(n6420), .ZN(n6295) );
  AOI22D0BWP U8512 ( .A1(n6466), .A2(N1105), .B1(n6467), .B2(N264), .ZN(n6420)
         );
  AOI221D0BWP U8513 ( .A1(vectorData2[32]), .A2(n6300), .B1(vectorData2[48]), 
        .B2(n6301), .C(n6469), .ZN(n6462) );
  AO22D0BWP U8514 ( .A1(n6303), .A2(vectorData2[240]), .B1(n6304), .B2(
        vectorData2[224]), .Z(n6469) );
  AO22D0BWP U8515 ( .A1(n6466), .A2(N1107), .B1(n6467), .B2(N266), .Z(n6304)
         );
  AO22D0BWP U8516 ( .A1(n6466), .A2(N1108), .B1(n6467), .B2(N267), .Z(n6303)
         );
  CKND0BWP U8517 ( .I(n6418), .ZN(n6301) );
  AOI22D0BWP U8518 ( .A1(n6466), .A2(N1096), .B1(n6467), .B2(N255), .ZN(n6418)
         );
  CKND0BWP U8519 ( .I(n6417), .ZN(n6300) );
  AOI22D0BWP U8520 ( .A1(n6466), .A2(N1095), .B1(n6467), .B2(N254), .ZN(n6417)
         );
  AOI222D0BWP U8521 ( .A1(vectorData2[96]), .A2(n6305), .B1(vectorData2[64]), 
        .B2(n6306), .C1(vectorData2[80]), .C2(n6307), .ZN(n6461) );
  CKND0BWP U8522 ( .I(n6414), .ZN(n6307) );
  AOI22D0BWP U8523 ( .A1(n6466), .A2(N1098), .B1(n6467), .B2(N257), .ZN(n6414)
         );
  CKND0BWP U8524 ( .I(n6415), .ZN(n6306) );
  AOI22D0BWP U8525 ( .A1(n6466), .A2(N1097), .B1(n6467), .B2(N256), .ZN(n6415)
         );
  CKND0BWP U8526 ( .I(n6416), .ZN(n6305) );
  AOI22D0BWP U8527 ( .A1(n6466), .A2(N1099), .B1(n6467), .B2(N258), .ZN(n6416)
         );
  OAI21D0BWP U8528 ( .A1(n6396), .A2(n6395), .B(n6404), .ZN(n6432) );
  IAO21D0BWP U8529 ( .A1(n6395), .A2(n5525), .B(n6344), .ZN(n6404) );
  INR2D0BWP U8530 ( .A1(n6470), .B1(n6395), .ZN(n6344) );
  ND3D0BWP U8531 ( .A1(code[1]), .A2(n6471), .A3(code[2]), .ZN(n5525) );
  CKND0BWP U8532 ( .I(n6409), .ZN(n6281) );
  NR2D0BWP U8533 ( .A1(n6406), .A2(n6395), .ZN(n6409) );
  CKND0BWP U8534 ( .I(n6285), .ZN(n6346) );
  NR2D0BWP U8535 ( .A1(n6472), .A2(n6395), .ZN(n6285) );
  NR2D0BWP U8536 ( .A1(n3368), .A2(n6209), .ZN(n6395) );
  OAI211D0BWP U8537 ( .A1(n6473), .A2(n6474), .B(n6475), .C(n6476), .ZN(N4085)
         );
  AOI222D0BWP U8538 ( .A1(Addr[15]), .A2(n6477), .B1(vectorData1[15]), .B2(
        n6478), .C1(scalarData1[15]), .C2(n6479), .ZN(n6476) );
  AOI22D0BWP U8539 ( .A1(n6480), .A2(n6481), .B1(n6482), .B2(n6483), .ZN(n6475) );
  ND4D0BWP U8540 ( .A1(n6484), .A2(n6485), .A3(n6486), .A4(n6487), .ZN(n6483)
         );
  AOI221D0BWP U8541 ( .A1(N1774), .A2(vectorData1[63]), .B1(N1775), .B2(
        vectorData1[79]), .C(n6488), .ZN(n6487) );
  OAI22D0BWP U8542 ( .A1(n6489), .A2(n6490), .B1(n6491), .B2(n6492), .ZN(n6488) );
  AOI221D0BWP U8543 ( .A1(N1778), .A2(vectorData1[127]), .B1(N1779), .B2(
        vectorData1[143]), .C(n6493), .ZN(n6486) );
  OAI22D0BWP U8544 ( .A1(n6494), .A2(n6495), .B1(n6496), .B2(n6497), .ZN(n6493) );
  AOI221D0BWP U8545 ( .A1(N1782), .A2(vectorData1[191]), .B1(N1783), .B2(
        vectorData1[207]), .C(n6498), .ZN(n6485) );
  OAI22D0BWP U8546 ( .A1(n6499), .A2(n6500), .B1(n6501), .B2(n6502), .ZN(n6498) );
  AOI222D0BWP U8547 ( .A1(N1786), .A2(vectorData1[255]), .B1(N1784), .B2(
        vectorData1[223]), .C1(N1785), .C2(vectorData1[239]), .ZN(n6484) );
  ND4D0BWP U8548 ( .A1(n6503), .A2(n6504), .A3(n6505), .A4(n6506), .ZN(n6481)
         );
  AOI221D0BWP U8549 ( .A1(vectorData1[63]), .A2(N255), .B1(vectorData1[79]), 
        .B2(N256), .C(n6507), .ZN(n6506) );
  OAI22D0BWP U8550 ( .A1(n6508), .A2(n6489), .B1(n6509), .B2(n6491), .ZN(n6507) );
  CKND0BWP U8551 ( .I(vectorData1[31]), .ZN(n6491) );
  CKND0BWP U8552 ( .I(vectorData1[47]), .ZN(n6489) );
  AOI221D0BWP U8553 ( .A1(vectorData1[127]), .A2(N259), .B1(vectorData1[143]), 
        .B2(N260), .C(n6510), .ZN(n6505) );
  OAI22D0BWP U8554 ( .A1(n6511), .A2(n6494), .B1(n6512), .B2(n6496), .ZN(n6510) );
  CKND0BWP U8555 ( .I(vectorData1[95]), .ZN(n6496) );
  CKND0BWP U8556 ( .I(vectorData1[111]), .ZN(n6494) );
  AOI221D0BWP U8557 ( .A1(vectorData1[191]), .A2(N263), .B1(vectorData1[207]), 
        .B2(N264), .C(n6513), .ZN(n6504) );
  OAI22D0BWP U8558 ( .A1(n6514), .A2(n6499), .B1(n6515), .B2(n6501), .ZN(n6513) );
  CKND0BWP U8559 ( .I(vectorData1[159]), .ZN(n6501) );
  CKND0BWP U8560 ( .I(vectorData1[175]), .ZN(n6499) );
  AOI222D0BWP U8561 ( .A1(vectorData1[255]), .A2(N267), .B1(vectorData1[223]), 
        .B2(N265), .C1(vectorData1[239]), .C2(N266), .ZN(n6503) );
  NR4D0BWP U8562 ( .A1(n6516), .A2(n6517), .A3(n6518), .A4(n6519), .ZN(n6473)
         );
  AO222D0BWP U8563 ( .A1(N1107), .A2(vectorData1[239]), .B1(N1106), .B2(
        vectorData1[223]), .C1(N1108), .C2(vectorData1[255]), .Z(n6519) );
  AO221D0BWP U8564 ( .A1(N1104), .A2(vectorData1[191]), .B1(N1105), .B2(
        vectorData1[207]), .C(n6520), .Z(n6518) );
  AO22D0BWP U8565 ( .A1(vectorData1[159]), .A2(N1102), .B1(vectorData1[175]), 
        .B2(N1103), .Z(n6520) );
  AO221D0BWP U8566 ( .A1(N1100), .A2(vectorData1[127]), .B1(N1101), .B2(
        vectorData1[143]), .C(n6521), .Z(n6517) );
  AO22D0BWP U8567 ( .A1(vectorData1[95]), .A2(N1098), .B1(vectorData1[111]), 
        .B2(N1099), .Z(n6521) );
  AO221D0BWP U8568 ( .A1(N1096), .A2(vectorData1[63]), .B1(N1097), .B2(
        vectorData1[79]), .C(n6522), .Z(n6516) );
  AO22D0BWP U8569 ( .A1(vectorData1[31]), .A2(N1094), .B1(vectorData1[47]), 
        .B2(N1095), .Z(n6522) );
  OAI211D0BWP U8570 ( .A1(n6523), .A2(n6474), .B(n6524), .C(n6525), .ZN(N4084)
         );
  AOI222D0BWP U8571 ( .A1(Addr[14]), .A2(n6477), .B1(vectorData1[14]), .B2(
        n6478), .C1(scalarData1[14]), .C2(n6479), .ZN(n6525) );
  AOI22D0BWP U8572 ( .A1(n6480), .A2(n6526), .B1(n6482), .B2(n6527), .ZN(n6524) );
  ND4D0BWP U8573 ( .A1(n6528), .A2(n6529), .A3(n6530), .A4(n6531), .ZN(n6527)
         );
  AOI221D0BWP U8574 ( .A1(vectorData1[62]), .A2(N1774), .B1(vectorData1[78]), 
        .B2(N1775), .C(n6532), .ZN(n6531) );
  OAI22D0BWP U8575 ( .A1(n6490), .A2(n6533), .B1(n6492), .B2(n6534), .ZN(n6532) );
  AOI221D0BWP U8576 ( .A1(vectorData1[126]), .A2(N1778), .B1(vectorData1[142]), 
        .B2(N1779), .C(n6535), .ZN(n6530) );
  OAI22D0BWP U8577 ( .A1(n6495), .A2(n6536), .B1(n6497), .B2(n6537), .ZN(n6535) );
  AOI221D0BWP U8578 ( .A1(vectorData1[190]), .A2(N1782), .B1(vectorData1[206]), 
        .B2(N1783), .C(n6538), .ZN(n6529) );
  OAI22D0BWP U8579 ( .A1(n6500), .A2(n6539), .B1(n6502), .B2(n6540), .ZN(n6538) );
  AOI222D0BWP U8580 ( .A1(vectorData1[254]), .A2(N1786), .B1(vectorData1[222]), 
        .B2(N1784), .C1(vectorData1[238]), .C2(N1785), .ZN(n6528) );
  ND4D0BWP U8581 ( .A1(n6541), .A2(n6542), .A3(n6543), .A4(n6544), .ZN(n6526)
         );
  AOI221D0BWP U8582 ( .A1(vectorData1[62]), .A2(N255), .B1(vectorData1[78]), 
        .B2(N256), .C(n6545), .ZN(n6544) );
  OAI22D0BWP U8583 ( .A1(n6508), .A2(n6533), .B1(n6509), .B2(n6534), .ZN(n6545) );
  CKND0BWP U8584 ( .I(vectorData1[30]), .ZN(n6534) );
  CKND0BWP U8585 ( .I(vectorData1[46]), .ZN(n6533) );
  AOI221D0BWP U8586 ( .A1(vectorData1[126]), .A2(N259), .B1(vectorData1[142]), 
        .B2(N260), .C(n6546), .ZN(n6543) );
  OAI22D0BWP U8587 ( .A1(n6511), .A2(n6536), .B1(n6512), .B2(n6537), .ZN(n6546) );
  CKND0BWP U8588 ( .I(vectorData1[94]), .ZN(n6537) );
  CKND0BWP U8589 ( .I(vectorData1[110]), .ZN(n6536) );
  AOI221D0BWP U8590 ( .A1(vectorData1[190]), .A2(N263), .B1(vectorData1[206]), 
        .B2(N264), .C(n6547), .ZN(n6542) );
  OAI22D0BWP U8591 ( .A1(n6514), .A2(n6539), .B1(n6515), .B2(n6540), .ZN(n6547) );
  CKND0BWP U8592 ( .I(vectorData1[158]), .ZN(n6540) );
  CKND0BWP U8593 ( .I(vectorData1[174]), .ZN(n6539) );
  AOI222D0BWP U8594 ( .A1(vectorData1[254]), .A2(N267), .B1(vectorData1[222]), 
        .B2(N265), .C1(vectorData1[238]), .C2(N266), .ZN(n6541) );
  NR4D0BWP U8595 ( .A1(n6548), .A2(n6549), .A3(n6550), .A4(n6551), .ZN(n6523)
         );
  AO222D0BWP U8596 ( .A1(N1107), .A2(vectorData1[238]), .B1(N1106), .B2(
        vectorData1[222]), .C1(N1108), .C2(vectorData1[254]), .Z(n6551) );
  AO221D0BWP U8597 ( .A1(N1104), .A2(vectorData1[190]), .B1(N1105), .B2(
        vectorData1[206]), .C(n6552), .Z(n6550) );
  AO22D0BWP U8598 ( .A1(vectorData1[158]), .A2(N1102), .B1(vectorData1[174]), 
        .B2(N1103), .Z(n6552) );
  AO221D0BWP U8599 ( .A1(N1100), .A2(vectorData1[126]), .B1(N1101), .B2(
        vectorData1[142]), .C(n6553), .Z(n6549) );
  AO22D0BWP U8600 ( .A1(vectorData1[94]), .A2(N1098), .B1(vectorData1[110]), 
        .B2(N1099), .Z(n6553) );
  AO221D0BWP U8601 ( .A1(N1096), .A2(vectorData1[62]), .B1(N1097), .B2(
        vectorData1[78]), .C(n6554), .Z(n6548) );
  AO22D0BWP U8602 ( .A1(vectorData1[30]), .A2(N1094), .B1(vectorData1[46]), 
        .B2(N1095), .Z(n6554) );
  OAI211D0BWP U8603 ( .A1(n6555), .A2(n6474), .B(n6556), .C(n6557), .ZN(N4083)
         );
  AOI222D0BWP U8604 ( .A1(Addr[13]), .A2(n6477), .B1(vectorData1[13]), .B2(
        n6478), .C1(scalarData1[13]), .C2(n6479), .ZN(n6557) );
  AOI22D0BWP U8605 ( .A1(n6480), .A2(n6558), .B1(n6482), .B2(n6559), .ZN(n6556) );
  ND4D0BWP U8606 ( .A1(n6560), .A2(n6561), .A3(n6562), .A4(n6563), .ZN(n6559)
         );
  AOI221D0BWP U8607 ( .A1(vectorData1[61]), .A2(N1774), .B1(vectorData1[77]), 
        .B2(N1775), .C(n6564), .ZN(n6563) );
  OAI22D0BWP U8608 ( .A1(n6490), .A2(n6565), .B1(n6492), .B2(n6566), .ZN(n6564) );
  AOI221D0BWP U8609 ( .A1(vectorData1[125]), .A2(N1778), .B1(vectorData1[141]), 
        .B2(N1779), .C(n6567), .ZN(n6562) );
  OAI22D0BWP U8610 ( .A1(n6495), .A2(n6568), .B1(n6497), .B2(n6569), .ZN(n6567) );
  AOI221D0BWP U8611 ( .A1(vectorData1[189]), .A2(N1782), .B1(vectorData1[205]), 
        .B2(N1783), .C(n6570), .ZN(n6561) );
  OAI22D0BWP U8612 ( .A1(n6500), .A2(n6571), .B1(n6502), .B2(n6572), .ZN(n6570) );
  AOI222D0BWP U8613 ( .A1(vectorData1[253]), .A2(N1786), .B1(vectorData1[221]), 
        .B2(N1784), .C1(vectorData1[237]), .C2(N1785), .ZN(n6560) );
  ND4D0BWP U8614 ( .A1(n6573), .A2(n6574), .A3(n6575), .A4(n6576), .ZN(n6558)
         );
  AOI221D0BWP U8615 ( .A1(vectorData1[61]), .A2(N255), .B1(vectorData1[77]), 
        .B2(N256), .C(n6577), .ZN(n6576) );
  OAI22D0BWP U8616 ( .A1(n6508), .A2(n6565), .B1(n6509), .B2(n6566), .ZN(n6577) );
  CKND0BWP U8617 ( .I(vectorData1[29]), .ZN(n6566) );
  CKND0BWP U8618 ( .I(vectorData1[45]), .ZN(n6565) );
  AOI221D0BWP U8619 ( .A1(vectorData1[125]), .A2(N259), .B1(vectorData1[141]), 
        .B2(N260), .C(n6578), .ZN(n6575) );
  OAI22D0BWP U8620 ( .A1(n6511), .A2(n6568), .B1(n6512), .B2(n6569), .ZN(n6578) );
  CKND0BWP U8621 ( .I(vectorData1[93]), .ZN(n6569) );
  CKND0BWP U8622 ( .I(vectorData1[109]), .ZN(n6568) );
  AOI221D0BWP U8623 ( .A1(vectorData1[189]), .A2(N263), .B1(vectorData1[205]), 
        .B2(N264), .C(n6579), .ZN(n6574) );
  OAI22D0BWP U8624 ( .A1(n6514), .A2(n6571), .B1(n6515), .B2(n6572), .ZN(n6579) );
  CKND0BWP U8625 ( .I(vectorData1[157]), .ZN(n6572) );
  CKND0BWP U8626 ( .I(vectorData1[173]), .ZN(n6571) );
  AOI222D0BWP U8627 ( .A1(vectorData1[253]), .A2(N267), .B1(vectorData1[221]), 
        .B2(N265), .C1(vectorData1[237]), .C2(N266), .ZN(n6573) );
  NR4D0BWP U8628 ( .A1(n6580), .A2(n6581), .A3(n6582), .A4(n6583), .ZN(n6555)
         );
  AO222D0BWP U8629 ( .A1(N1107), .A2(vectorData1[237]), .B1(N1106), .B2(
        vectorData1[221]), .C1(N1108), .C2(vectorData1[253]), .Z(n6583) );
  AO221D0BWP U8630 ( .A1(N1104), .A2(vectorData1[189]), .B1(N1105), .B2(
        vectorData1[205]), .C(n6584), .Z(n6582) );
  AO22D0BWP U8631 ( .A1(vectorData1[157]), .A2(N1102), .B1(vectorData1[173]), 
        .B2(N1103), .Z(n6584) );
  AO221D0BWP U8632 ( .A1(N1100), .A2(vectorData1[125]), .B1(N1101), .B2(
        vectorData1[141]), .C(n6585), .Z(n6581) );
  AO22D0BWP U8633 ( .A1(vectorData1[93]), .A2(N1098), .B1(vectorData1[109]), 
        .B2(N1099), .Z(n6585) );
  AO221D0BWP U8634 ( .A1(N1096), .A2(vectorData1[61]), .B1(N1097), .B2(
        vectorData1[77]), .C(n6586), .Z(n6580) );
  AO22D0BWP U8635 ( .A1(vectorData1[29]), .A2(N1094), .B1(vectorData1[45]), 
        .B2(N1095), .Z(n6586) );
  OAI211D0BWP U8636 ( .A1(n6587), .A2(n6474), .B(n6588), .C(n6589), .ZN(N4082)
         );
  AOI222D0BWP U8637 ( .A1(Addr[12]), .A2(n6477), .B1(vectorData1[12]), .B2(
        n6478), .C1(scalarData1[12]), .C2(n6479), .ZN(n6589) );
  AOI22D0BWP U8638 ( .A1(n6480), .A2(n6590), .B1(n6482), .B2(n6591), .ZN(n6588) );
  ND4D0BWP U8639 ( .A1(n6592), .A2(n6593), .A3(n6594), .A4(n6595), .ZN(n6591)
         );
  AOI221D0BWP U8640 ( .A1(vectorData1[60]), .A2(N1774), .B1(vectorData1[76]), 
        .B2(N1775), .C(n6596), .ZN(n6595) );
  OAI22D0BWP U8641 ( .A1(n6490), .A2(n6597), .B1(n6492), .B2(n6598), .ZN(n6596) );
  AOI221D0BWP U8642 ( .A1(vectorData1[124]), .A2(N1778), .B1(vectorData1[140]), 
        .B2(N1779), .C(n6599), .ZN(n6594) );
  OAI22D0BWP U8643 ( .A1(n6495), .A2(n6600), .B1(n6497), .B2(n6601), .ZN(n6599) );
  AOI221D0BWP U8644 ( .A1(vectorData1[188]), .A2(N1782), .B1(vectorData1[204]), 
        .B2(N1783), .C(n6602), .ZN(n6593) );
  OAI22D0BWP U8645 ( .A1(n6500), .A2(n6603), .B1(n6502), .B2(n6604), .ZN(n6602) );
  AOI222D0BWP U8646 ( .A1(vectorData1[252]), .A2(N1786), .B1(vectorData1[220]), 
        .B2(N1784), .C1(vectorData1[236]), .C2(N1785), .ZN(n6592) );
  ND4D0BWP U8647 ( .A1(n6605), .A2(n6606), .A3(n6607), .A4(n6608), .ZN(n6590)
         );
  AOI221D0BWP U8648 ( .A1(vectorData1[60]), .A2(N255), .B1(vectorData1[76]), 
        .B2(N256), .C(n6609), .ZN(n6608) );
  OAI22D0BWP U8649 ( .A1(n6508), .A2(n6597), .B1(n6509), .B2(n6598), .ZN(n6609) );
  CKND0BWP U8650 ( .I(vectorData1[28]), .ZN(n6598) );
  CKND0BWP U8651 ( .I(vectorData1[44]), .ZN(n6597) );
  AOI221D0BWP U8652 ( .A1(vectorData1[124]), .A2(N259), .B1(vectorData1[140]), 
        .B2(N260), .C(n6610), .ZN(n6607) );
  OAI22D0BWP U8653 ( .A1(n6511), .A2(n6600), .B1(n6512), .B2(n6601), .ZN(n6610) );
  CKND0BWP U8654 ( .I(vectorData1[92]), .ZN(n6601) );
  CKND0BWP U8655 ( .I(vectorData1[108]), .ZN(n6600) );
  AOI221D0BWP U8656 ( .A1(vectorData1[188]), .A2(N263), .B1(vectorData1[204]), 
        .B2(N264), .C(n6611), .ZN(n6606) );
  OAI22D0BWP U8657 ( .A1(n6514), .A2(n6603), .B1(n6515), .B2(n6604), .ZN(n6611) );
  CKND0BWP U8658 ( .I(vectorData1[156]), .ZN(n6604) );
  CKND0BWP U8659 ( .I(vectorData1[172]), .ZN(n6603) );
  AOI222D0BWP U8660 ( .A1(vectorData1[252]), .A2(N267), .B1(vectorData1[220]), 
        .B2(N265), .C1(vectorData1[236]), .C2(N266), .ZN(n6605) );
  NR4D0BWP U8661 ( .A1(n6612), .A2(n6613), .A3(n6614), .A4(n6615), .ZN(n6587)
         );
  AO222D0BWP U8662 ( .A1(N1107), .A2(vectorData1[236]), .B1(N1106), .B2(
        vectorData1[220]), .C1(N1108), .C2(vectorData1[252]), .Z(n6615) );
  AO221D0BWP U8663 ( .A1(N1104), .A2(vectorData1[188]), .B1(N1105), .B2(
        vectorData1[204]), .C(n6616), .Z(n6614) );
  AO22D0BWP U8664 ( .A1(vectorData1[156]), .A2(N1102), .B1(vectorData1[172]), 
        .B2(N1103), .Z(n6616) );
  AO221D0BWP U8665 ( .A1(N1100), .A2(vectorData1[124]), .B1(N1101), .B2(
        vectorData1[140]), .C(n6617), .Z(n6613) );
  AO22D0BWP U8666 ( .A1(vectorData1[92]), .A2(N1098), .B1(vectorData1[108]), 
        .B2(N1099), .Z(n6617) );
  AO221D0BWP U8667 ( .A1(N1096), .A2(vectorData1[60]), .B1(N1097), .B2(
        vectorData1[76]), .C(n6618), .Z(n6612) );
  AO22D0BWP U8668 ( .A1(vectorData1[28]), .A2(N1094), .B1(vectorData1[44]), 
        .B2(N1095), .Z(n6618) );
  OAI211D0BWP U8669 ( .A1(n6619), .A2(n6474), .B(n6620), .C(n6621), .ZN(N4081)
         );
  AOI222D0BWP U8670 ( .A1(Addr[11]), .A2(n6477), .B1(vectorData1[11]), .B2(
        n6478), .C1(scalarData1[11]), .C2(n6479), .ZN(n6621) );
  AOI22D0BWP U8671 ( .A1(n6480), .A2(n6622), .B1(n6482), .B2(n6623), .ZN(n6620) );
  ND4D0BWP U8672 ( .A1(n6624), .A2(n6625), .A3(n6626), .A4(n6627), .ZN(n6623)
         );
  AOI221D0BWP U8673 ( .A1(vectorData1[59]), .A2(N1774), .B1(vectorData1[75]), 
        .B2(N1775), .C(n6628), .ZN(n6627) );
  OAI22D0BWP U8674 ( .A1(n6490), .A2(n6629), .B1(n6492), .B2(n6630), .ZN(n6628) );
  AOI221D0BWP U8675 ( .A1(vectorData1[123]), .A2(N1778), .B1(vectorData1[139]), 
        .B2(N1779), .C(n6631), .ZN(n6626) );
  OAI22D0BWP U8676 ( .A1(n6495), .A2(n6632), .B1(n6497), .B2(n6633), .ZN(n6631) );
  AOI221D0BWP U8677 ( .A1(vectorData1[187]), .A2(N1782), .B1(vectorData1[203]), 
        .B2(N1783), .C(n6634), .ZN(n6625) );
  OAI22D0BWP U8678 ( .A1(n6500), .A2(n6635), .B1(n6502), .B2(n6636), .ZN(n6634) );
  AOI222D0BWP U8679 ( .A1(vectorData1[251]), .A2(N1786), .B1(vectorData1[219]), 
        .B2(N1784), .C1(vectorData1[235]), .C2(N1785), .ZN(n6624) );
  ND4D0BWP U8680 ( .A1(n6637), .A2(n6638), .A3(n6639), .A4(n6640), .ZN(n6622)
         );
  AOI221D0BWP U8681 ( .A1(vectorData1[59]), .A2(N255), .B1(vectorData1[75]), 
        .B2(N256), .C(n6641), .ZN(n6640) );
  OAI22D0BWP U8682 ( .A1(n6508), .A2(n6629), .B1(n6509), .B2(n6630), .ZN(n6641) );
  CKND0BWP U8683 ( .I(vectorData1[27]), .ZN(n6630) );
  CKND0BWP U8684 ( .I(vectorData1[43]), .ZN(n6629) );
  AOI221D0BWP U8685 ( .A1(vectorData1[123]), .A2(N259), .B1(vectorData1[139]), 
        .B2(N260), .C(n6642), .ZN(n6639) );
  OAI22D0BWP U8686 ( .A1(n6511), .A2(n6632), .B1(n6512), .B2(n6633), .ZN(n6642) );
  CKND0BWP U8687 ( .I(vectorData1[91]), .ZN(n6633) );
  CKND0BWP U8688 ( .I(vectorData1[107]), .ZN(n6632) );
  AOI221D0BWP U8689 ( .A1(vectorData1[187]), .A2(N263), .B1(vectorData1[203]), 
        .B2(N264), .C(n6643), .ZN(n6638) );
  OAI22D0BWP U8690 ( .A1(n6514), .A2(n6635), .B1(n6515), .B2(n6636), .ZN(n6643) );
  CKND0BWP U8691 ( .I(vectorData1[155]), .ZN(n6636) );
  CKND0BWP U8692 ( .I(vectorData1[171]), .ZN(n6635) );
  AOI222D0BWP U8693 ( .A1(vectorData1[251]), .A2(N267), .B1(vectorData1[219]), 
        .B2(N265), .C1(vectorData1[235]), .C2(N266), .ZN(n6637) );
  NR4D0BWP U8694 ( .A1(n6644), .A2(n6645), .A3(n6646), .A4(n6647), .ZN(n6619)
         );
  AO222D0BWP U8695 ( .A1(N1107), .A2(vectorData1[235]), .B1(N1106), .B2(
        vectorData1[219]), .C1(N1108), .C2(vectorData1[251]), .Z(n6647) );
  AO221D0BWP U8696 ( .A1(N1104), .A2(vectorData1[187]), .B1(N1105), .B2(
        vectorData1[203]), .C(n6648), .Z(n6646) );
  AO22D0BWP U8697 ( .A1(vectorData1[155]), .A2(N1102), .B1(vectorData1[171]), 
        .B2(N1103), .Z(n6648) );
  AO221D0BWP U8698 ( .A1(N1100), .A2(vectorData1[123]), .B1(N1101), .B2(
        vectorData1[139]), .C(n6649), .Z(n6645) );
  AO22D0BWP U8699 ( .A1(vectorData1[91]), .A2(N1098), .B1(vectorData1[107]), 
        .B2(N1099), .Z(n6649) );
  AO221D0BWP U8700 ( .A1(N1096), .A2(vectorData1[59]), .B1(N1097), .B2(
        vectorData1[75]), .C(n6650), .Z(n6644) );
  AO22D0BWP U8701 ( .A1(vectorData1[27]), .A2(N1094), .B1(vectorData1[43]), 
        .B2(N1095), .Z(n6650) );
  OAI211D0BWP U8702 ( .A1(n6651), .A2(n6474), .B(n6652), .C(n6653), .ZN(N4080)
         );
  AOI222D0BWP U8703 ( .A1(Addr[10]), .A2(n6477), .B1(vectorData1[10]), .B2(
        n6478), .C1(scalarData1[10]), .C2(n6479), .ZN(n6653) );
  AOI22D0BWP U8704 ( .A1(n6480), .A2(n6654), .B1(n6482), .B2(n6655), .ZN(n6652) );
  ND4D0BWP U8705 ( .A1(n6656), .A2(n6657), .A3(n6658), .A4(n6659), .ZN(n6655)
         );
  AOI221D0BWP U8706 ( .A1(vectorData1[58]), .A2(N1774), .B1(vectorData1[74]), 
        .B2(N1775), .C(n6660), .ZN(n6659) );
  OAI22D0BWP U8707 ( .A1(n6490), .A2(n6661), .B1(n6492), .B2(n6662), .ZN(n6660) );
  AOI221D0BWP U8708 ( .A1(vectorData1[122]), .A2(N1778), .B1(vectorData1[138]), 
        .B2(N1779), .C(n6663), .ZN(n6658) );
  OAI22D0BWP U8709 ( .A1(n6495), .A2(n6664), .B1(n6497), .B2(n6665), .ZN(n6663) );
  AOI221D0BWP U8710 ( .A1(vectorData1[186]), .A2(N1782), .B1(vectorData1[202]), 
        .B2(N1783), .C(n6666), .ZN(n6657) );
  OAI22D0BWP U8711 ( .A1(n6500), .A2(n6667), .B1(n6502), .B2(n6668), .ZN(n6666) );
  AOI222D0BWP U8712 ( .A1(vectorData1[250]), .A2(N1786), .B1(vectorData1[218]), 
        .B2(N1784), .C1(vectorData1[234]), .C2(N1785), .ZN(n6656) );
  ND4D0BWP U8713 ( .A1(n6669), .A2(n6670), .A3(n6671), .A4(n6672), .ZN(n6654)
         );
  AOI221D0BWP U8714 ( .A1(vectorData1[58]), .A2(N255), .B1(vectorData1[74]), 
        .B2(N256), .C(n6673), .ZN(n6672) );
  OAI22D0BWP U8715 ( .A1(n6508), .A2(n6661), .B1(n6509), .B2(n6662), .ZN(n6673) );
  CKND0BWP U8716 ( .I(vectorData1[26]), .ZN(n6662) );
  CKND0BWP U8717 ( .I(vectorData1[42]), .ZN(n6661) );
  AOI221D0BWP U8718 ( .A1(vectorData1[122]), .A2(N259), .B1(vectorData1[138]), 
        .B2(N260), .C(n6674), .ZN(n6671) );
  OAI22D0BWP U8719 ( .A1(n6511), .A2(n6664), .B1(n6512), .B2(n6665), .ZN(n6674) );
  CKND0BWP U8720 ( .I(vectorData1[90]), .ZN(n6665) );
  CKND0BWP U8721 ( .I(vectorData1[106]), .ZN(n6664) );
  AOI221D0BWP U8722 ( .A1(vectorData1[186]), .A2(N263), .B1(vectorData1[202]), 
        .B2(N264), .C(n6675), .ZN(n6670) );
  OAI22D0BWP U8723 ( .A1(n6514), .A2(n6667), .B1(n6515), .B2(n6668), .ZN(n6675) );
  CKND0BWP U8724 ( .I(vectorData1[154]), .ZN(n6668) );
  CKND0BWP U8725 ( .I(vectorData1[170]), .ZN(n6667) );
  AOI222D0BWP U8726 ( .A1(vectorData1[250]), .A2(N267), .B1(vectorData1[218]), 
        .B2(N265), .C1(vectorData1[234]), .C2(N266), .ZN(n6669) );
  NR4D0BWP U8727 ( .A1(n6676), .A2(n6677), .A3(n6678), .A4(n6679), .ZN(n6651)
         );
  AO222D0BWP U8728 ( .A1(N1107), .A2(vectorData1[234]), .B1(N1106), .B2(
        vectorData1[218]), .C1(N1108), .C2(vectorData1[250]), .Z(n6679) );
  AO221D0BWP U8729 ( .A1(N1104), .A2(vectorData1[186]), .B1(N1105), .B2(
        vectorData1[202]), .C(n6680), .Z(n6678) );
  AO22D0BWP U8730 ( .A1(vectorData1[154]), .A2(N1102), .B1(vectorData1[170]), 
        .B2(N1103), .Z(n6680) );
  AO221D0BWP U8731 ( .A1(N1100), .A2(vectorData1[122]), .B1(N1101), .B2(
        vectorData1[138]), .C(n6681), .Z(n6677) );
  AO22D0BWP U8732 ( .A1(vectorData1[90]), .A2(N1098), .B1(vectorData1[106]), 
        .B2(N1099), .Z(n6681) );
  AO221D0BWP U8733 ( .A1(N1096), .A2(vectorData1[58]), .B1(N1097), .B2(
        vectorData1[74]), .C(n6682), .Z(n6676) );
  AO22D0BWP U8734 ( .A1(vectorData1[26]), .A2(N1094), .B1(vectorData1[42]), 
        .B2(N1095), .Z(n6682) );
  OAI211D0BWP U8735 ( .A1(n6683), .A2(n6474), .B(n6684), .C(n6685), .ZN(N4079)
         );
  AOI222D0BWP U8736 ( .A1(Addr[9]), .A2(n6477), .B1(vectorData1[9]), .B2(n6478), .C1(scalarData1[9]), .C2(n6479), .ZN(n6685) );
  AOI22D0BWP U8737 ( .A1(n6480), .A2(n6686), .B1(n6482), .B2(n6687), .ZN(n6684) );
  ND4D0BWP U8738 ( .A1(n6688), .A2(n6689), .A3(n6690), .A4(n6691), .ZN(n6687)
         );
  AOI221D0BWP U8739 ( .A1(vectorData1[57]), .A2(N1774), .B1(vectorData1[73]), 
        .B2(N1775), .C(n6692), .ZN(n6691) );
  OAI22D0BWP U8740 ( .A1(n6490), .A2(n6693), .B1(n6492), .B2(n6694), .ZN(n6692) );
  AOI221D0BWP U8741 ( .A1(vectorData1[121]), .A2(N1778), .B1(vectorData1[137]), 
        .B2(N1779), .C(n6695), .ZN(n6690) );
  OAI22D0BWP U8742 ( .A1(n6495), .A2(n6696), .B1(n6497), .B2(n6697), .ZN(n6695) );
  AOI221D0BWP U8743 ( .A1(vectorData1[185]), .A2(N1782), .B1(vectorData1[201]), 
        .B2(N1783), .C(n6698), .ZN(n6689) );
  OAI22D0BWP U8744 ( .A1(n6500), .A2(n6699), .B1(n6502), .B2(n6700), .ZN(n6698) );
  AOI222D0BWP U8745 ( .A1(vectorData1[249]), .A2(N1786), .B1(vectorData1[217]), 
        .B2(N1784), .C1(vectorData1[233]), .C2(N1785), .ZN(n6688) );
  ND4D0BWP U8746 ( .A1(n6701), .A2(n6702), .A3(n6703), .A4(n6704), .ZN(n6686)
         );
  AOI221D0BWP U8747 ( .A1(vectorData1[57]), .A2(N255), .B1(vectorData1[73]), 
        .B2(N256), .C(n6705), .ZN(n6704) );
  OAI22D0BWP U8748 ( .A1(n6508), .A2(n6693), .B1(n6509), .B2(n6694), .ZN(n6705) );
  CKND0BWP U8749 ( .I(vectorData1[25]), .ZN(n6694) );
  CKND0BWP U8750 ( .I(vectorData1[41]), .ZN(n6693) );
  AOI221D0BWP U8751 ( .A1(vectorData1[121]), .A2(N259), .B1(vectorData1[137]), 
        .B2(N260), .C(n6706), .ZN(n6703) );
  OAI22D0BWP U8752 ( .A1(n6511), .A2(n6696), .B1(n6512), .B2(n6697), .ZN(n6706) );
  CKND0BWP U8753 ( .I(vectorData1[89]), .ZN(n6697) );
  CKND0BWP U8754 ( .I(vectorData1[105]), .ZN(n6696) );
  AOI221D0BWP U8755 ( .A1(vectorData1[185]), .A2(N263), .B1(vectorData1[201]), 
        .B2(N264), .C(n6707), .ZN(n6702) );
  OAI22D0BWP U8756 ( .A1(n6514), .A2(n6699), .B1(n6515), .B2(n6700), .ZN(n6707) );
  CKND0BWP U8757 ( .I(vectorData1[153]), .ZN(n6700) );
  CKND0BWP U8758 ( .I(vectorData1[169]), .ZN(n6699) );
  AOI222D0BWP U8759 ( .A1(vectorData1[249]), .A2(N267), .B1(vectorData1[217]), 
        .B2(N265), .C1(vectorData1[233]), .C2(N266), .ZN(n6701) );
  NR4D0BWP U8760 ( .A1(n6708), .A2(n6709), .A3(n6710), .A4(n6711), .ZN(n6683)
         );
  AO222D0BWP U8761 ( .A1(N1107), .A2(vectorData1[233]), .B1(N1106), .B2(
        vectorData1[217]), .C1(N1108), .C2(vectorData1[249]), .Z(n6711) );
  AO221D0BWP U8762 ( .A1(N1104), .A2(vectorData1[185]), .B1(N1105), .B2(
        vectorData1[201]), .C(n6712), .Z(n6710) );
  AO22D0BWP U8763 ( .A1(vectorData1[153]), .A2(N1102), .B1(vectorData1[169]), 
        .B2(N1103), .Z(n6712) );
  AO221D0BWP U8764 ( .A1(N1100), .A2(vectorData1[121]), .B1(N1101), .B2(
        vectorData1[137]), .C(n6713), .Z(n6709) );
  AO22D0BWP U8765 ( .A1(vectorData1[89]), .A2(N1098), .B1(vectorData1[105]), 
        .B2(N1099), .Z(n6713) );
  AO221D0BWP U8766 ( .A1(N1096), .A2(vectorData1[57]), .B1(N1097), .B2(
        vectorData1[73]), .C(n6714), .Z(n6708) );
  AO22D0BWP U8767 ( .A1(vectorData1[25]), .A2(N1094), .B1(vectorData1[41]), 
        .B2(N1095), .Z(n6714) );
  OAI211D0BWP U8768 ( .A1(n6715), .A2(n6474), .B(n6716), .C(n6717), .ZN(N4078)
         );
  AOI222D0BWP U8769 ( .A1(Addr[8]), .A2(n6477), .B1(vectorData1[8]), .B2(n6478), .C1(scalarData1[8]), .C2(n6479), .ZN(n6717) );
  AOI22D0BWP U8770 ( .A1(n6480), .A2(n6718), .B1(n6482), .B2(n6719), .ZN(n6716) );
  ND4D0BWP U8771 ( .A1(n6720), .A2(n6721), .A3(n6722), .A4(n6723), .ZN(n6719)
         );
  AOI221D0BWP U8772 ( .A1(vectorData1[56]), .A2(N1774), .B1(vectorData1[72]), 
        .B2(N1775), .C(n6724), .ZN(n6723) );
  OAI22D0BWP U8773 ( .A1(n6490), .A2(n6725), .B1(n6492), .B2(n6726), .ZN(n6724) );
  AOI221D0BWP U8774 ( .A1(vectorData1[120]), .A2(N1778), .B1(vectorData1[136]), 
        .B2(N1779), .C(n6727), .ZN(n6722) );
  OAI22D0BWP U8775 ( .A1(n6495), .A2(n6728), .B1(n6497), .B2(n6729), .ZN(n6727) );
  AOI221D0BWP U8776 ( .A1(vectorData1[184]), .A2(N1782), .B1(vectorData1[200]), 
        .B2(N1783), .C(n6730), .ZN(n6721) );
  OAI22D0BWP U8777 ( .A1(n6500), .A2(n6731), .B1(n6502), .B2(n6732), .ZN(n6730) );
  AOI222D0BWP U8778 ( .A1(vectorData1[248]), .A2(N1786), .B1(vectorData1[216]), 
        .B2(N1784), .C1(vectorData1[232]), .C2(N1785), .ZN(n6720) );
  ND4D0BWP U8779 ( .A1(n6733), .A2(n6734), .A3(n6735), .A4(n6736), .ZN(n6718)
         );
  AOI221D0BWP U8780 ( .A1(vectorData1[56]), .A2(N255), .B1(vectorData1[72]), 
        .B2(N256), .C(n6737), .ZN(n6736) );
  OAI22D0BWP U8781 ( .A1(n6508), .A2(n6725), .B1(n6509), .B2(n6726), .ZN(n6737) );
  CKND0BWP U8782 ( .I(vectorData1[24]), .ZN(n6726) );
  CKND0BWP U8783 ( .I(vectorData1[40]), .ZN(n6725) );
  AOI221D0BWP U8784 ( .A1(vectorData1[120]), .A2(N259), .B1(vectorData1[136]), 
        .B2(N260), .C(n6738), .ZN(n6735) );
  OAI22D0BWP U8785 ( .A1(n6511), .A2(n6728), .B1(n6512), .B2(n6729), .ZN(n6738) );
  CKND0BWP U8786 ( .I(vectorData1[88]), .ZN(n6729) );
  CKND0BWP U8787 ( .I(vectorData1[104]), .ZN(n6728) );
  AOI221D0BWP U8788 ( .A1(vectorData1[184]), .A2(N263), .B1(vectorData1[200]), 
        .B2(N264), .C(n6739), .ZN(n6734) );
  OAI22D0BWP U8789 ( .A1(n6514), .A2(n6731), .B1(n6515), .B2(n6732), .ZN(n6739) );
  CKND0BWP U8790 ( .I(vectorData1[152]), .ZN(n6732) );
  CKND0BWP U8791 ( .I(vectorData1[168]), .ZN(n6731) );
  AOI222D0BWP U8792 ( .A1(vectorData1[248]), .A2(N267), .B1(vectorData1[216]), 
        .B2(N265), .C1(vectorData1[232]), .C2(N266), .ZN(n6733) );
  NR4D0BWP U8793 ( .A1(n6740), .A2(n6741), .A3(n6742), .A4(n6743), .ZN(n6715)
         );
  AO222D0BWP U8794 ( .A1(N1107), .A2(vectorData1[232]), .B1(N1106), .B2(
        vectorData1[216]), .C1(N1108), .C2(vectorData1[248]), .Z(n6743) );
  AO221D0BWP U8795 ( .A1(N1104), .A2(vectorData1[184]), .B1(N1105), .B2(
        vectorData1[200]), .C(n6744), .Z(n6742) );
  AO22D0BWP U8796 ( .A1(vectorData1[152]), .A2(N1102), .B1(vectorData1[168]), 
        .B2(N1103), .Z(n6744) );
  AO221D0BWP U8797 ( .A1(N1100), .A2(vectorData1[120]), .B1(N1101), .B2(
        vectorData1[136]), .C(n6745), .Z(n6741) );
  AO22D0BWP U8798 ( .A1(vectorData1[88]), .A2(N1098), .B1(vectorData1[104]), 
        .B2(N1099), .Z(n6745) );
  AO221D0BWP U8799 ( .A1(N1096), .A2(vectorData1[56]), .B1(N1097), .B2(
        vectorData1[72]), .C(n6746), .Z(n6740) );
  AO22D0BWP U8800 ( .A1(vectorData1[24]), .A2(N1094), .B1(vectorData1[40]), 
        .B2(N1095), .Z(n6746) );
  OAI211D0BWP U8801 ( .A1(n6747), .A2(n6474), .B(n6748), .C(n6749), .ZN(N4077)
         );
  AOI222D0BWP U8802 ( .A1(Addr[7]), .A2(n6477), .B1(vectorData1[7]), .B2(n6478), .C1(scalarData1[7]), .C2(n6479), .ZN(n6749) );
  AOI22D0BWP U8803 ( .A1(n6480), .A2(n6750), .B1(n6482), .B2(n6751), .ZN(n6748) );
  ND4D0BWP U8804 ( .A1(n6752), .A2(n6753), .A3(n6754), .A4(n6755), .ZN(n6751)
         );
  AOI221D0BWP U8805 ( .A1(vectorData1[55]), .A2(N1774), .B1(vectorData1[71]), 
        .B2(N1775), .C(n6756), .ZN(n6755) );
  OAI22D0BWP U8806 ( .A1(n6490), .A2(n6757), .B1(n6492), .B2(n6758), .ZN(n6756) );
  AOI221D0BWP U8807 ( .A1(vectorData1[119]), .A2(N1778), .B1(vectorData1[135]), 
        .B2(N1779), .C(n6759), .ZN(n6754) );
  OAI22D0BWP U8808 ( .A1(n6495), .A2(n6760), .B1(n6497), .B2(n6761), .ZN(n6759) );
  AOI221D0BWP U8809 ( .A1(vectorData1[183]), .A2(N1782), .B1(vectorData1[199]), 
        .B2(N1783), .C(n6762), .ZN(n6753) );
  OAI22D0BWP U8810 ( .A1(n6500), .A2(n6763), .B1(n6502), .B2(n6764), .ZN(n6762) );
  AOI222D0BWP U8811 ( .A1(vectorData1[247]), .A2(N1786), .B1(vectorData1[215]), 
        .B2(N1784), .C1(vectorData1[231]), .C2(N1785), .ZN(n6752) );
  ND4D0BWP U8812 ( .A1(n6765), .A2(n6766), .A3(n6767), .A4(n6768), .ZN(n6750)
         );
  AOI221D0BWP U8813 ( .A1(vectorData1[55]), .A2(N255), .B1(vectorData1[71]), 
        .B2(N256), .C(n6769), .ZN(n6768) );
  OAI22D0BWP U8814 ( .A1(n6508), .A2(n6757), .B1(n6509), .B2(n6758), .ZN(n6769) );
  CKND0BWP U8815 ( .I(vectorData1[23]), .ZN(n6758) );
  CKND0BWP U8816 ( .I(vectorData1[39]), .ZN(n6757) );
  AOI221D0BWP U8817 ( .A1(vectorData1[119]), .A2(N259), .B1(vectorData1[135]), 
        .B2(N260), .C(n6770), .ZN(n6767) );
  OAI22D0BWP U8818 ( .A1(n6511), .A2(n6760), .B1(n6512), .B2(n6761), .ZN(n6770) );
  CKND0BWP U8819 ( .I(vectorData1[87]), .ZN(n6761) );
  CKND0BWP U8820 ( .I(vectorData1[103]), .ZN(n6760) );
  AOI221D0BWP U8821 ( .A1(vectorData1[183]), .A2(N263), .B1(vectorData1[199]), 
        .B2(N264), .C(n6771), .ZN(n6766) );
  OAI22D0BWP U8822 ( .A1(n6514), .A2(n6763), .B1(n6515), .B2(n6764), .ZN(n6771) );
  CKND0BWP U8823 ( .I(vectorData1[151]), .ZN(n6764) );
  CKND0BWP U8824 ( .I(vectorData1[167]), .ZN(n6763) );
  AOI222D0BWP U8825 ( .A1(vectorData1[247]), .A2(N267), .B1(vectorData1[215]), 
        .B2(N265), .C1(vectorData1[231]), .C2(N266), .ZN(n6765) );
  NR4D0BWP U8826 ( .A1(n6772), .A2(n6773), .A3(n6774), .A4(n6775), .ZN(n6747)
         );
  AO222D0BWP U8827 ( .A1(N1107), .A2(vectorData1[231]), .B1(N1106), .B2(
        vectorData1[215]), .C1(N1108), .C2(vectorData1[247]), .Z(n6775) );
  AO221D0BWP U8828 ( .A1(N1104), .A2(vectorData1[183]), .B1(N1105), .B2(
        vectorData1[199]), .C(n6776), .Z(n6774) );
  AO22D0BWP U8829 ( .A1(vectorData1[151]), .A2(N1102), .B1(vectorData1[167]), 
        .B2(N1103), .Z(n6776) );
  AO221D0BWP U8830 ( .A1(N1100), .A2(vectorData1[119]), .B1(N1101), .B2(
        vectorData1[135]), .C(n6777), .Z(n6773) );
  AO22D0BWP U8831 ( .A1(vectorData1[87]), .A2(N1098), .B1(vectorData1[103]), 
        .B2(N1099), .Z(n6777) );
  AO221D0BWP U8832 ( .A1(N1096), .A2(vectorData1[55]), .B1(N1097), .B2(
        vectorData1[71]), .C(n6778), .Z(n6772) );
  AO22D0BWP U8833 ( .A1(vectorData1[23]), .A2(N1094), .B1(vectorData1[39]), 
        .B2(N1095), .Z(n6778) );
  OAI211D0BWP U8834 ( .A1(n6779), .A2(n6474), .B(n6780), .C(n6781), .ZN(N4076)
         );
  AOI222D0BWP U8835 ( .A1(Addr[6]), .A2(n6477), .B1(vectorData1[6]), .B2(n6478), .C1(scalarData1[6]), .C2(n6479), .ZN(n6781) );
  AOI22D0BWP U8836 ( .A1(n6480), .A2(n6782), .B1(n6482), .B2(n6783), .ZN(n6780) );
  ND4D0BWP U8837 ( .A1(n6784), .A2(n6785), .A3(n6786), .A4(n6787), .ZN(n6783)
         );
  AOI221D0BWP U8838 ( .A1(vectorData1[54]), .A2(N1774), .B1(vectorData1[70]), 
        .B2(N1775), .C(n6788), .ZN(n6787) );
  OAI22D0BWP U8839 ( .A1(n6490), .A2(n6789), .B1(n6492), .B2(n6790), .ZN(n6788) );
  AOI221D0BWP U8840 ( .A1(vectorData1[118]), .A2(N1778), .B1(vectorData1[134]), 
        .B2(N1779), .C(n6791), .ZN(n6786) );
  OAI22D0BWP U8841 ( .A1(n6495), .A2(n6792), .B1(n6497), .B2(n6793), .ZN(n6791) );
  AOI221D0BWP U8842 ( .A1(vectorData1[182]), .A2(N1782), .B1(vectorData1[198]), 
        .B2(N1783), .C(n6794), .ZN(n6785) );
  OAI22D0BWP U8843 ( .A1(n6500), .A2(n6795), .B1(n6502), .B2(n6796), .ZN(n6794) );
  AOI222D0BWP U8844 ( .A1(vectorData1[246]), .A2(N1786), .B1(vectorData1[214]), 
        .B2(N1784), .C1(vectorData1[230]), .C2(N1785), .ZN(n6784) );
  ND4D0BWP U8845 ( .A1(n6797), .A2(n6798), .A3(n6799), .A4(n6800), .ZN(n6782)
         );
  AOI221D0BWP U8846 ( .A1(vectorData1[54]), .A2(N255), .B1(vectorData1[70]), 
        .B2(N256), .C(n6801), .ZN(n6800) );
  OAI22D0BWP U8847 ( .A1(n6508), .A2(n6789), .B1(n6509), .B2(n6790), .ZN(n6801) );
  CKND0BWP U8848 ( .I(vectorData1[22]), .ZN(n6790) );
  CKND0BWP U8849 ( .I(vectorData1[38]), .ZN(n6789) );
  AOI221D0BWP U8850 ( .A1(vectorData1[118]), .A2(N259), .B1(vectorData1[134]), 
        .B2(N260), .C(n6802), .ZN(n6799) );
  OAI22D0BWP U8851 ( .A1(n6511), .A2(n6792), .B1(n6512), .B2(n6793), .ZN(n6802) );
  CKND0BWP U8852 ( .I(vectorData1[86]), .ZN(n6793) );
  CKND0BWP U8853 ( .I(vectorData1[102]), .ZN(n6792) );
  AOI221D0BWP U8854 ( .A1(vectorData1[182]), .A2(N263), .B1(vectorData1[198]), 
        .B2(N264), .C(n6803), .ZN(n6798) );
  OAI22D0BWP U8855 ( .A1(n6514), .A2(n6795), .B1(n6515), .B2(n6796), .ZN(n6803) );
  CKND0BWP U8856 ( .I(vectorData1[150]), .ZN(n6796) );
  CKND0BWP U8857 ( .I(vectorData1[166]), .ZN(n6795) );
  AOI222D0BWP U8858 ( .A1(vectorData1[246]), .A2(N267), .B1(vectorData1[214]), 
        .B2(N265), .C1(vectorData1[230]), .C2(N266), .ZN(n6797) );
  NR4D0BWP U8859 ( .A1(n6804), .A2(n6805), .A3(n6806), .A4(n6807), .ZN(n6779)
         );
  AO222D0BWP U8860 ( .A1(N1107), .A2(vectorData1[230]), .B1(N1106), .B2(
        vectorData1[214]), .C1(N1108), .C2(vectorData1[246]), .Z(n6807) );
  AO221D0BWP U8861 ( .A1(N1104), .A2(vectorData1[182]), .B1(N1105), .B2(
        vectorData1[198]), .C(n6808), .Z(n6806) );
  AO22D0BWP U8862 ( .A1(vectorData1[150]), .A2(N1102), .B1(vectorData1[166]), 
        .B2(N1103), .Z(n6808) );
  AO221D0BWP U8863 ( .A1(N1100), .A2(vectorData1[118]), .B1(N1101), .B2(
        vectorData1[134]), .C(n6809), .Z(n6805) );
  AO22D0BWP U8864 ( .A1(vectorData1[86]), .A2(N1098), .B1(vectorData1[102]), 
        .B2(N1099), .Z(n6809) );
  AO221D0BWP U8865 ( .A1(N1096), .A2(vectorData1[54]), .B1(N1097), .B2(
        vectorData1[70]), .C(n6810), .Z(n6804) );
  AO22D0BWP U8866 ( .A1(vectorData1[22]), .A2(N1094), .B1(vectorData1[38]), 
        .B2(N1095), .Z(n6810) );
  OAI211D0BWP U8867 ( .A1(n6811), .A2(n6474), .B(n6812), .C(n6813), .ZN(N4075)
         );
  AOI222D0BWP U8868 ( .A1(Addr[5]), .A2(n6477), .B1(vectorData1[5]), .B2(n6478), .C1(scalarData1[5]), .C2(n6479), .ZN(n6813) );
  AOI22D0BWP U8869 ( .A1(n6480), .A2(n6814), .B1(n6482), .B2(n6815), .ZN(n6812) );
  ND4D0BWP U8870 ( .A1(n6816), .A2(n6817), .A3(n6818), .A4(n6819), .ZN(n6815)
         );
  AOI221D0BWP U8871 ( .A1(vectorData1[53]), .A2(N1774), .B1(vectorData1[69]), 
        .B2(N1775), .C(n6820), .ZN(n6819) );
  OAI22D0BWP U8872 ( .A1(n6490), .A2(n6821), .B1(n6492), .B2(n6822), .ZN(n6820) );
  AOI221D0BWP U8873 ( .A1(vectorData1[117]), .A2(N1778), .B1(vectorData1[133]), 
        .B2(N1779), .C(n6823), .ZN(n6818) );
  OAI22D0BWP U8874 ( .A1(n6495), .A2(n6824), .B1(n6497), .B2(n6825), .ZN(n6823) );
  AOI221D0BWP U8875 ( .A1(vectorData1[181]), .A2(N1782), .B1(vectorData1[197]), 
        .B2(N1783), .C(n6826), .ZN(n6817) );
  OAI22D0BWP U8876 ( .A1(n6500), .A2(n6827), .B1(n6502), .B2(n6828), .ZN(n6826) );
  AOI222D0BWP U8877 ( .A1(vectorData1[245]), .A2(N1786), .B1(vectorData1[213]), 
        .B2(N1784), .C1(vectorData1[229]), .C2(N1785), .ZN(n6816) );
  ND4D0BWP U8878 ( .A1(n6829), .A2(n6830), .A3(n6831), .A4(n6832), .ZN(n6814)
         );
  AOI221D0BWP U8879 ( .A1(vectorData1[53]), .A2(N255), .B1(vectorData1[69]), 
        .B2(N256), .C(n6833), .ZN(n6832) );
  OAI22D0BWP U8880 ( .A1(n6508), .A2(n6821), .B1(n6509), .B2(n6822), .ZN(n6833) );
  CKND0BWP U8881 ( .I(vectorData1[21]), .ZN(n6822) );
  CKND0BWP U8882 ( .I(vectorData1[37]), .ZN(n6821) );
  AOI221D0BWP U8883 ( .A1(vectorData1[117]), .A2(N259), .B1(vectorData1[133]), 
        .B2(N260), .C(n6834), .ZN(n6831) );
  OAI22D0BWP U8884 ( .A1(n6511), .A2(n6824), .B1(n6512), .B2(n6825), .ZN(n6834) );
  CKND0BWP U8885 ( .I(vectorData1[85]), .ZN(n6825) );
  CKND0BWP U8886 ( .I(vectorData1[101]), .ZN(n6824) );
  AOI221D0BWP U8887 ( .A1(vectorData1[181]), .A2(N263), .B1(vectorData1[197]), 
        .B2(N264), .C(n6835), .ZN(n6830) );
  OAI22D0BWP U8888 ( .A1(n6514), .A2(n6827), .B1(n6515), .B2(n6828), .ZN(n6835) );
  CKND0BWP U8889 ( .I(vectorData1[149]), .ZN(n6828) );
  CKND0BWP U8890 ( .I(vectorData1[165]), .ZN(n6827) );
  AOI222D0BWP U8891 ( .A1(vectorData1[245]), .A2(N267), .B1(vectorData1[213]), 
        .B2(N265), .C1(vectorData1[229]), .C2(N266), .ZN(n6829) );
  NR4D0BWP U8892 ( .A1(n6836), .A2(n6837), .A3(n6838), .A4(n6839), .ZN(n6811)
         );
  AO222D0BWP U8893 ( .A1(N1107), .A2(vectorData1[229]), .B1(N1106), .B2(
        vectorData1[213]), .C1(N1108), .C2(vectorData1[245]), .Z(n6839) );
  AO221D0BWP U8894 ( .A1(N1104), .A2(vectorData1[181]), .B1(N1105), .B2(
        vectorData1[197]), .C(n6840), .Z(n6838) );
  AO22D0BWP U8895 ( .A1(vectorData1[149]), .A2(N1102), .B1(vectorData1[165]), 
        .B2(N1103), .Z(n6840) );
  AO221D0BWP U8896 ( .A1(N1100), .A2(vectorData1[117]), .B1(N1101), .B2(
        vectorData1[133]), .C(n6841), .Z(n6837) );
  AO22D0BWP U8897 ( .A1(vectorData1[85]), .A2(N1098), .B1(vectorData1[101]), 
        .B2(N1099), .Z(n6841) );
  AO221D0BWP U8898 ( .A1(N1096), .A2(vectorData1[53]), .B1(N1097), .B2(
        vectorData1[69]), .C(n6842), .Z(n6836) );
  AO22D0BWP U8899 ( .A1(vectorData1[21]), .A2(N1094), .B1(vectorData1[37]), 
        .B2(N1095), .Z(n6842) );
  OAI211D0BWP U8900 ( .A1(n6843), .A2(n6474), .B(n6844), .C(n6845), .ZN(N4074)
         );
  AOI222D0BWP U8901 ( .A1(Addr[4]), .A2(n6477), .B1(vectorData1[4]), .B2(n6478), .C1(scalarData1[4]), .C2(n6479), .ZN(n6845) );
  AOI22D0BWP U8902 ( .A1(n6480), .A2(n6846), .B1(n6482), .B2(n6847), .ZN(n6844) );
  ND4D0BWP U8903 ( .A1(n6848), .A2(n6849), .A3(n6850), .A4(n6851), .ZN(n6847)
         );
  AOI221D0BWP U8904 ( .A1(vectorData1[52]), .A2(N1774), .B1(vectorData1[68]), 
        .B2(N1775), .C(n6852), .ZN(n6851) );
  OAI22D0BWP U8905 ( .A1(n6490), .A2(n6853), .B1(n6492), .B2(n6854), .ZN(n6852) );
  AOI221D0BWP U8906 ( .A1(vectorData1[116]), .A2(N1778), .B1(vectorData1[132]), 
        .B2(N1779), .C(n6855), .ZN(n6850) );
  OAI22D0BWP U8907 ( .A1(n6495), .A2(n6856), .B1(n6497), .B2(n6857), .ZN(n6855) );
  AOI221D0BWP U8908 ( .A1(vectorData1[180]), .A2(N1782), .B1(vectorData1[196]), 
        .B2(N1783), .C(n6858), .ZN(n6849) );
  OAI22D0BWP U8909 ( .A1(n6500), .A2(n6859), .B1(n6502), .B2(n6860), .ZN(n6858) );
  AOI222D0BWP U8910 ( .A1(vectorData1[244]), .A2(N1786), .B1(vectorData1[212]), 
        .B2(N1784), .C1(vectorData1[228]), .C2(N1785), .ZN(n6848) );
  ND4D0BWP U8911 ( .A1(n6861), .A2(n6862), .A3(n6863), .A4(n6864), .ZN(n6846)
         );
  AOI221D0BWP U8912 ( .A1(vectorData1[52]), .A2(N255), .B1(vectorData1[68]), 
        .B2(N256), .C(n6865), .ZN(n6864) );
  OAI22D0BWP U8913 ( .A1(n6508), .A2(n6853), .B1(n6509), .B2(n6854), .ZN(n6865) );
  CKND0BWP U8914 ( .I(vectorData1[20]), .ZN(n6854) );
  CKND0BWP U8915 ( .I(vectorData1[36]), .ZN(n6853) );
  AOI221D0BWP U8916 ( .A1(vectorData1[116]), .A2(N259), .B1(vectorData1[132]), 
        .B2(N260), .C(n6866), .ZN(n6863) );
  OAI22D0BWP U8917 ( .A1(n6511), .A2(n6856), .B1(n6512), .B2(n6857), .ZN(n6866) );
  CKND0BWP U8918 ( .I(vectorData1[84]), .ZN(n6857) );
  CKND0BWP U8919 ( .I(vectorData1[100]), .ZN(n6856) );
  AOI221D0BWP U8920 ( .A1(vectorData1[180]), .A2(N263), .B1(vectorData1[196]), 
        .B2(N264), .C(n6867), .ZN(n6862) );
  OAI22D0BWP U8921 ( .A1(n6514), .A2(n6859), .B1(n6515), .B2(n6860), .ZN(n6867) );
  CKND0BWP U8922 ( .I(vectorData1[148]), .ZN(n6860) );
  CKND0BWP U8923 ( .I(vectorData1[164]), .ZN(n6859) );
  AOI222D0BWP U8924 ( .A1(vectorData1[244]), .A2(N267), .B1(vectorData1[212]), 
        .B2(N265), .C1(vectorData1[228]), .C2(N266), .ZN(n6861) );
  NR4D0BWP U8925 ( .A1(n6868), .A2(n6869), .A3(n6870), .A4(n6871), .ZN(n6843)
         );
  AO222D0BWP U8926 ( .A1(N1107), .A2(vectorData1[228]), .B1(N1106), .B2(
        vectorData1[212]), .C1(N1108), .C2(vectorData1[244]), .Z(n6871) );
  AO221D0BWP U8927 ( .A1(N1104), .A2(vectorData1[180]), .B1(N1105), .B2(
        vectorData1[196]), .C(n6872), .Z(n6870) );
  AO22D0BWP U8928 ( .A1(vectorData1[148]), .A2(N1102), .B1(vectorData1[164]), 
        .B2(N1103), .Z(n6872) );
  AO221D0BWP U8929 ( .A1(N1100), .A2(vectorData1[116]), .B1(N1101), .B2(
        vectorData1[132]), .C(n6873), .Z(n6869) );
  AO22D0BWP U8930 ( .A1(vectorData1[84]), .A2(N1098), .B1(vectorData1[100]), 
        .B2(N1099), .Z(n6873) );
  AO221D0BWP U8931 ( .A1(N1096), .A2(vectorData1[52]), .B1(N1097), .B2(
        vectorData1[68]), .C(n6874), .Z(n6868) );
  AO22D0BWP U8932 ( .A1(vectorData1[20]), .A2(N1094), .B1(vectorData1[36]), 
        .B2(N1095), .Z(n6874) );
  OAI211D0BWP U8933 ( .A1(n6875), .A2(n6474), .B(n6876), .C(n6877), .ZN(N4073)
         );
  AOI222D0BWP U8934 ( .A1(Addr[3]), .A2(n6477), .B1(vectorData1[3]), .B2(n6478), .C1(scalarData1[3]), .C2(n6479), .ZN(n6877) );
  AOI22D0BWP U8935 ( .A1(n6480), .A2(n6878), .B1(n6482), .B2(n6879), .ZN(n6876) );
  ND4D0BWP U8936 ( .A1(n6880), .A2(n6881), .A3(n6882), .A4(n6883), .ZN(n6879)
         );
  AOI221D0BWP U8937 ( .A1(vectorData1[51]), .A2(N1774), .B1(vectorData1[67]), 
        .B2(N1775), .C(n6884), .ZN(n6883) );
  OAI22D0BWP U8938 ( .A1(n6490), .A2(n6885), .B1(n6492), .B2(n6886), .ZN(n6884) );
  AOI221D0BWP U8939 ( .A1(vectorData1[115]), .A2(N1778), .B1(vectorData1[131]), 
        .B2(N1779), .C(n6887), .ZN(n6882) );
  OAI22D0BWP U8940 ( .A1(n6495), .A2(n6888), .B1(n6497), .B2(n6889), .ZN(n6887) );
  AOI221D0BWP U8941 ( .A1(vectorData1[179]), .A2(N1782), .B1(vectorData1[195]), 
        .B2(N1783), .C(n6890), .ZN(n6881) );
  OAI22D0BWP U8942 ( .A1(n6500), .A2(n6891), .B1(n6502), .B2(n6892), .ZN(n6890) );
  AOI222D0BWP U8943 ( .A1(vectorData1[243]), .A2(N1786), .B1(vectorData1[211]), 
        .B2(N1784), .C1(vectorData1[227]), .C2(N1785), .ZN(n6880) );
  ND4D0BWP U8944 ( .A1(n6893), .A2(n6894), .A3(n6895), .A4(n6896), .ZN(n6878)
         );
  AOI221D0BWP U8945 ( .A1(vectorData1[51]), .A2(N255), .B1(vectorData1[67]), 
        .B2(N256), .C(n6897), .ZN(n6896) );
  OAI22D0BWP U8946 ( .A1(n6508), .A2(n6885), .B1(n6509), .B2(n6886), .ZN(n6897) );
  CKND0BWP U8947 ( .I(vectorData1[19]), .ZN(n6886) );
  CKND0BWP U8948 ( .I(vectorData1[35]), .ZN(n6885) );
  AOI221D0BWP U8949 ( .A1(vectorData1[115]), .A2(N259), .B1(vectorData1[131]), 
        .B2(N260), .C(n6898), .ZN(n6895) );
  OAI22D0BWP U8950 ( .A1(n6511), .A2(n6888), .B1(n6512), .B2(n6889), .ZN(n6898) );
  CKND0BWP U8951 ( .I(vectorData1[83]), .ZN(n6889) );
  CKND0BWP U8952 ( .I(vectorData1[99]), .ZN(n6888) );
  AOI221D0BWP U8953 ( .A1(vectorData1[179]), .A2(N263), .B1(vectorData1[195]), 
        .B2(N264), .C(n6899), .ZN(n6894) );
  OAI22D0BWP U8954 ( .A1(n6514), .A2(n6891), .B1(n6515), .B2(n6892), .ZN(n6899) );
  CKND0BWP U8955 ( .I(vectorData1[147]), .ZN(n6892) );
  CKND0BWP U8956 ( .I(vectorData1[163]), .ZN(n6891) );
  AOI222D0BWP U8957 ( .A1(vectorData1[243]), .A2(N267), .B1(vectorData1[211]), 
        .B2(N265), .C1(vectorData1[227]), .C2(N266), .ZN(n6893) );
  NR4D0BWP U8958 ( .A1(n6900), .A2(n6901), .A3(n6902), .A4(n6903), .ZN(n6875)
         );
  AO222D0BWP U8959 ( .A1(N1107), .A2(vectorData1[227]), .B1(N1106), .B2(
        vectorData1[211]), .C1(N1108), .C2(vectorData1[243]), .Z(n6903) );
  AO221D0BWP U8960 ( .A1(N1104), .A2(vectorData1[179]), .B1(N1105), .B2(
        vectorData1[195]), .C(n6904), .Z(n6902) );
  AO22D0BWP U8961 ( .A1(vectorData1[147]), .A2(N1102), .B1(vectorData1[163]), 
        .B2(N1103), .Z(n6904) );
  AO221D0BWP U8962 ( .A1(N1100), .A2(vectorData1[115]), .B1(N1101), .B2(
        vectorData1[131]), .C(n6905), .Z(n6901) );
  AO22D0BWP U8963 ( .A1(vectorData1[83]), .A2(N1098), .B1(vectorData1[99]), 
        .B2(N1099), .Z(n6905) );
  AO221D0BWP U8964 ( .A1(N1096), .A2(vectorData1[51]), .B1(N1097), .B2(
        vectorData1[67]), .C(n6906), .Z(n6900) );
  AO22D0BWP U8965 ( .A1(vectorData1[19]), .A2(N1094), .B1(vectorData1[35]), 
        .B2(N1095), .Z(n6906) );
  OAI211D0BWP U8966 ( .A1(n6907), .A2(n6474), .B(n6908), .C(n6909), .ZN(N4072)
         );
  AOI222D0BWP U8967 ( .A1(Addr[2]), .A2(n6477), .B1(vectorData1[2]), .B2(n6478), .C1(scalarData1[2]), .C2(n6479), .ZN(n6909) );
  AOI22D0BWP U8968 ( .A1(n6480), .A2(n6910), .B1(n6482), .B2(n6911), .ZN(n6908) );
  ND4D0BWP U8969 ( .A1(n6912), .A2(n6913), .A3(n6914), .A4(n6915), .ZN(n6911)
         );
  AOI221D0BWP U8970 ( .A1(vectorData1[50]), .A2(N1774), .B1(vectorData1[66]), 
        .B2(N1775), .C(n6916), .ZN(n6915) );
  OAI22D0BWP U8971 ( .A1(n6490), .A2(n6917), .B1(n6492), .B2(n6918), .ZN(n6916) );
  AOI221D0BWP U8972 ( .A1(vectorData1[114]), .A2(N1778), .B1(vectorData1[130]), 
        .B2(N1779), .C(n6919), .ZN(n6914) );
  OAI22D0BWP U8973 ( .A1(n6495), .A2(n6920), .B1(n6497), .B2(n6921), .ZN(n6919) );
  AOI221D0BWP U8974 ( .A1(vectorData1[178]), .A2(N1782), .B1(vectorData1[194]), 
        .B2(N1783), .C(n6922), .ZN(n6913) );
  OAI22D0BWP U8975 ( .A1(n6500), .A2(n6923), .B1(n6502), .B2(n6924), .ZN(n6922) );
  AOI222D0BWP U8976 ( .A1(vectorData1[242]), .A2(N1786), .B1(vectorData1[210]), 
        .B2(N1784), .C1(vectorData1[226]), .C2(N1785), .ZN(n6912) );
  ND4D0BWP U8977 ( .A1(n6925), .A2(n6926), .A3(n6927), .A4(n6928), .ZN(n6910)
         );
  AOI221D0BWP U8978 ( .A1(vectorData1[50]), .A2(N255), .B1(vectorData1[66]), 
        .B2(N256), .C(n6929), .ZN(n6928) );
  OAI22D0BWP U8979 ( .A1(n6508), .A2(n6917), .B1(n6509), .B2(n6918), .ZN(n6929) );
  CKND0BWP U8980 ( .I(vectorData1[18]), .ZN(n6918) );
  CKND0BWP U8981 ( .I(vectorData1[34]), .ZN(n6917) );
  AOI221D0BWP U8982 ( .A1(vectorData1[114]), .A2(N259), .B1(vectorData1[130]), 
        .B2(N260), .C(n6930), .ZN(n6927) );
  OAI22D0BWP U8983 ( .A1(n6511), .A2(n6920), .B1(n6512), .B2(n6921), .ZN(n6930) );
  CKND0BWP U8984 ( .I(vectorData1[82]), .ZN(n6921) );
  CKND0BWP U8985 ( .I(vectorData1[98]), .ZN(n6920) );
  AOI221D0BWP U8986 ( .A1(vectorData1[178]), .A2(N263), .B1(vectorData1[194]), 
        .B2(N264), .C(n6931), .ZN(n6926) );
  OAI22D0BWP U8987 ( .A1(n6514), .A2(n6923), .B1(n6515), .B2(n6924), .ZN(n6931) );
  CKND0BWP U8988 ( .I(vectorData1[146]), .ZN(n6924) );
  CKND0BWP U8989 ( .I(vectorData1[162]), .ZN(n6923) );
  AOI222D0BWP U8990 ( .A1(vectorData1[242]), .A2(N267), .B1(vectorData1[210]), 
        .B2(N265), .C1(vectorData1[226]), .C2(N266), .ZN(n6925) );
  NR4D0BWP U8991 ( .A1(n6932), .A2(n6933), .A3(n6934), .A4(n6935), .ZN(n6907)
         );
  AO222D0BWP U8992 ( .A1(N1107), .A2(vectorData1[226]), .B1(N1106), .B2(
        vectorData1[210]), .C1(N1108), .C2(vectorData1[242]), .Z(n6935) );
  AO221D0BWP U8993 ( .A1(N1104), .A2(vectorData1[178]), .B1(N1105), .B2(
        vectorData1[194]), .C(n6936), .Z(n6934) );
  AO22D0BWP U8994 ( .A1(vectorData1[146]), .A2(N1102), .B1(vectorData1[162]), 
        .B2(N1103), .Z(n6936) );
  AO221D0BWP U8995 ( .A1(N1100), .A2(vectorData1[114]), .B1(N1101), .B2(
        vectorData1[130]), .C(n6937), .Z(n6933) );
  AO22D0BWP U8996 ( .A1(vectorData1[82]), .A2(N1098), .B1(vectorData1[98]), 
        .B2(N1099), .Z(n6937) );
  AO221D0BWP U8997 ( .A1(N1096), .A2(vectorData1[50]), .B1(N1097), .B2(
        vectorData1[66]), .C(n6938), .Z(n6932) );
  AO22D0BWP U8998 ( .A1(vectorData1[18]), .A2(N1094), .B1(vectorData1[34]), 
        .B2(N1095), .Z(n6938) );
  OAI211D0BWP U8999 ( .A1(n6939), .A2(n6474), .B(n6940), .C(n6941), .ZN(N4071)
         );
  AOI222D0BWP U9000 ( .A1(Addr[1]), .A2(n6477), .B1(vectorData1[1]), .B2(n6478), .C1(scalarData1[1]), .C2(n6479), .ZN(n6941) );
  AOI22D0BWP U9001 ( .A1(n6480), .A2(n6942), .B1(n6482), .B2(n6943), .ZN(n6940) );
  ND4D0BWP U9002 ( .A1(n6944), .A2(n6945), .A3(n6946), .A4(n6947), .ZN(n6943)
         );
  AOI221D0BWP U9003 ( .A1(vectorData1[49]), .A2(N1774), .B1(vectorData1[65]), 
        .B2(N1775), .C(n6948), .ZN(n6947) );
  OAI22D0BWP U9004 ( .A1(n6490), .A2(n6949), .B1(n6492), .B2(n6950), .ZN(n6948) );
  AOI221D0BWP U9005 ( .A1(vectorData1[113]), .A2(N1778), .B1(vectorData1[129]), 
        .B2(N1779), .C(n6951), .ZN(n6946) );
  OAI22D0BWP U9006 ( .A1(n6495), .A2(n6952), .B1(n6497), .B2(n6953), .ZN(n6951) );
  AOI221D0BWP U9007 ( .A1(vectorData1[177]), .A2(N1782), .B1(vectorData1[193]), 
        .B2(N1783), .C(n6954), .ZN(n6945) );
  OAI22D0BWP U9008 ( .A1(n6500), .A2(n6955), .B1(n6502), .B2(n6956), .ZN(n6954) );
  AOI222D0BWP U9009 ( .A1(vectorData1[241]), .A2(N1786), .B1(vectorData1[209]), 
        .B2(N1784), .C1(vectorData1[225]), .C2(N1785), .ZN(n6944) );
  ND4D0BWP U9010 ( .A1(n6957), .A2(n6958), .A3(n6959), .A4(n6960), .ZN(n6942)
         );
  AOI221D0BWP U9011 ( .A1(vectorData1[49]), .A2(N255), .B1(vectorData1[65]), 
        .B2(N256), .C(n6961), .ZN(n6960) );
  OAI22D0BWP U9012 ( .A1(n6508), .A2(n6949), .B1(n6509), .B2(n6950), .ZN(n6961) );
  CKND0BWP U9013 ( .I(vectorData1[17]), .ZN(n6950) );
  CKND0BWP U9014 ( .I(vectorData1[33]), .ZN(n6949) );
  AOI221D0BWP U9015 ( .A1(vectorData1[113]), .A2(N259), .B1(vectorData1[129]), 
        .B2(N260), .C(n6962), .ZN(n6959) );
  OAI22D0BWP U9016 ( .A1(n6511), .A2(n6952), .B1(n6512), .B2(n6953), .ZN(n6962) );
  CKND0BWP U9017 ( .I(vectorData1[81]), .ZN(n6953) );
  CKND0BWP U9018 ( .I(vectorData1[97]), .ZN(n6952) );
  AOI221D0BWP U9019 ( .A1(vectorData1[177]), .A2(N263), .B1(vectorData1[193]), 
        .B2(N264), .C(n6963), .ZN(n6958) );
  OAI22D0BWP U9020 ( .A1(n6514), .A2(n6955), .B1(n6515), .B2(n6956), .ZN(n6963) );
  CKND0BWP U9021 ( .I(vectorData1[145]), .ZN(n6956) );
  CKND0BWP U9022 ( .I(vectorData1[161]), .ZN(n6955) );
  AOI222D0BWP U9023 ( .A1(vectorData1[241]), .A2(N267), .B1(vectorData1[209]), 
        .B2(N265), .C1(vectorData1[225]), .C2(N266), .ZN(n6957) );
  NR4D0BWP U9024 ( .A1(n6964), .A2(n6965), .A3(n6966), .A4(n6967), .ZN(n6939)
         );
  AO222D0BWP U9025 ( .A1(N1107), .A2(vectorData1[225]), .B1(N1106), .B2(
        vectorData1[209]), .C1(N1108), .C2(vectorData1[241]), .Z(n6967) );
  AO221D0BWP U9026 ( .A1(N1104), .A2(vectorData1[177]), .B1(N1105), .B2(
        vectorData1[193]), .C(n6968), .Z(n6966) );
  AO22D0BWP U9027 ( .A1(vectorData1[145]), .A2(N1102), .B1(vectorData1[161]), 
        .B2(N1103), .Z(n6968) );
  AO221D0BWP U9028 ( .A1(N1100), .A2(vectorData1[113]), .B1(N1101), .B2(
        vectorData1[129]), .C(n6969), .Z(n6965) );
  AO22D0BWP U9029 ( .A1(vectorData1[81]), .A2(N1098), .B1(vectorData1[97]), 
        .B2(N1099), .Z(n6969) );
  AO221D0BWP U9030 ( .A1(N1096), .A2(vectorData1[49]), .B1(N1097), .B2(
        vectorData1[65]), .C(n6970), .Z(n6964) );
  AO22D0BWP U9031 ( .A1(vectorData1[17]), .A2(N1094), .B1(vectorData1[33]), 
        .B2(N1095), .Z(n6970) );
  OAI211D0BWP U9032 ( .A1(n6971), .A2(n6474), .B(n6972), .C(n6973), .ZN(N4070)
         );
  AOI222D0BWP U9033 ( .A1(Addr[0]), .A2(n6477), .B1(vectorData1[0]), .B2(n6478), .C1(scalarData1[0]), .C2(n6479), .ZN(n6973) );
  OA211D0BWP U9034 ( .A1(n6974), .A2(code[2]), .B(n6471), .C(n3368), .Z(n6479)
         );
  NR2D0BWP U9035 ( .A1(n6198), .A2(n6975), .ZN(n6974) );
  INR2D0BWP U9036 ( .A1(n6976), .B1(n6250), .ZN(n6478) );
  CKND0BWP U9037 ( .I(n6977), .ZN(n6477) );
  AOI22D0BWP U9038 ( .A1(n6480), .A2(n6978), .B1(n6482), .B2(n6979), .ZN(n6972) );
  ND4D0BWP U9039 ( .A1(n6980), .A2(n6981), .A3(n6982), .A4(n6983), .ZN(n6979)
         );
  AOI221D0BWP U9040 ( .A1(vectorData1[48]), .A2(N1774), .B1(vectorData1[64]), 
        .B2(N1775), .C(n6984), .ZN(n6983) );
  OAI22D0BWP U9041 ( .A1(n6490), .A2(n6985), .B1(n6492), .B2(n6986), .ZN(n6984) );
  CKND0BWP U9042 ( .I(N1772), .ZN(n6492) );
  CKND0BWP U9043 ( .I(N1773), .ZN(n6490) );
  AOI221D0BWP U9044 ( .A1(vectorData1[112]), .A2(N1778), .B1(vectorData1[128]), 
        .B2(N1779), .C(n6987), .ZN(n6982) );
  OAI22D0BWP U9045 ( .A1(n6495), .A2(n6988), .B1(n6497), .B2(n6989), .ZN(n6987) );
  CKND0BWP U9046 ( .I(N1776), .ZN(n6497) );
  CKND0BWP U9047 ( .I(N1777), .ZN(n6495) );
  AOI221D0BWP U9048 ( .A1(vectorData1[176]), .A2(N1782), .B1(vectorData1[192]), 
        .B2(N1783), .C(n6990), .ZN(n6981) );
  OAI22D0BWP U9049 ( .A1(n6500), .A2(n6991), .B1(n6502), .B2(n6992), .ZN(n6990) );
  CKND0BWP U9050 ( .I(N1780), .ZN(n6502) );
  CKND0BWP U9051 ( .I(N1781), .ZN(n6500) );
  AOI222D0BWP U9052 ( .A1(vectorData1[240]), .A2(N1786), .B1(vectorData1[208]), 
        .B2(N1784), .C1(vectorData1[224]), .C2(N1785), .ZN(n6980) );
  INR2D0BWP U9053 ( .A1(n6976), .B1(n6993), .ZN(n6482) );
  ND4D0BWP U9054 ( .A1(n6994), .A2(n6995), .A3(n6996), .A4(n6997), .ZN(n6978)
         );
  AOI221D0BWP U9055 ( .A1(vectorData1[48]), .A2(N255), .B1(vectorData1[64]), 
        .B2(N256), .C(n6998), .ZN(n6997) );
  OAI22D0BWP U9056 ( .A1(n6508), .A2(n6985), .B1(n6509), .B2(n6986), .ZN(n6998) );
  CKND0BWP U9057 ( .I(vectorData1[16]), .ZN(n6986) );
  CKND0BWP U9058 ( .I(N253), .ZN(n6509) );
  CKND0BWP U9059 ( .I(vectorData1[32]), .ZN(n6985) );
  CKND0BWP U9060 ( .I(N254), .ZN(n6508) );
  AOI221D0BWP U9061 ( .A1(vectorData1[112]), .A2(N259), .B1(vectorData1[128]), 
        .B2(N260), .C(n6999), .ZN(n6996) );
  OAI22D0BWP U9062 ( .A1(n6511), .A2(n6988), .B1(n6512), .B2(n6989), .ZN(n6999) );
  CKND0BWP U9063 ( .I(vectorData1[80]), .ZN(n6989) );
  CKND0BWP U9064 ( .I(N257), .ZN(n6512) );
  CKND0BWP U9065 ( .I(vectorData1[96]), .ZN(n6988) );
  CKND0BWP U9066 ( .I(N258), .ZN(n6511) );
  AOI221D0BWP U9067 ( .A1(vectorData1[176]), .A2(N263), .B1(vectorData1[192]), 
        .B2(N264), .C(n7000), .ZN(n6995) );
  OAI22D0BWP U9068 ( .A1(n6514), .A2(n6991), .B1(n6515), .B2(n6992), .ZN(n7000) );
  CKND0BWP U9069 ( .I(vectorData1[144]), .ZN(n6992) );
  CKND0BWP U9070 ( .I(N261), .ZN(n6515) );
  CKND0BWP U9071 ( .I(vectorData1[160]), .ZN(n6991) );
  CKND0BWP U9072 ( .I(N262), .ZN(n6514) );
  AOI222D0BWP U9073 ( .A1(vectorData1[240]), .A2(N267), .B1(vectorData1[208]), 
        .B2(N265), .C1(vectorData1[224]), .C2(N266), .ZN(n6994) );
  INR2D0BWP U9074 ( .A1(n6976), .B1(n6169), .ZN(n6480) );
  CKND2D0BWP U9075 ( .A1(n6976), .A2(n6466), .ZN(n6474) );
  CKND2D0BWP U9076 ( .A1(n6472), .A2(n6406), .ZN(n6976) );
  NR4D0BWP U9077 ( .A1(n7001), .A2(n7002), .A3(n7003), .A4(n7004), .ZN(n6971)
         );
  AO222D0BWP U9078 ( .A1(N1107), .A2(vectorData1[224]), .B1(N1106), .B2(
        vectorData1[208]), .C1(N1108), .C2(vectorData1[240]), .Z(n7004) );
  AO221D0BWP U9079 ( .A1(N1104), .A2(vectorData1[176]), .B1(N1105), .B2(
        vectorData1[192]), .C(n7005), .Z(n7003) );
  AO22D0BWP U9080 ( .A1(vectorData1[144]), .A2(N1102), .B1(vectorData1[160]), 
        .B2(N1103), .Z(n7005) );
  AO221D0BWP U9081 ( .A1(N1100), .A2(vectorData1[112]), .B1(N1101), .B2(
        vectorData1[128]), .C(n7006), .Z(n7002) );
  AO22D0BWP U9082 ( .A1(vectorData1[80]), .A2(N1098), .B1(vectorData1[96]), 
        .B2(N1099), .Z(n7006) );
  AO221D0BWP U9083 ( .A1(N1096), .A2(vectorData1[48]), .B1(N1097), .B2(
        vectorData1[64]), .C(n7007), .Z(n7001) );
  AO22D0BWP U9084 ( .A1(vectorData1[16]), .A2(N1094), .B1(vectorData1[32]), 
        .B2(N1095), .Z(n7007) );
  OAI22D0BWP U9085 ( .A1(n7008), .A2(n7009), .B1(n2522), .B2(n7010), .ZN(N4069) );
  AOI21D0BWP U9086 ( .A1(cycles[4]), .A2(n7011), .B(n5600), .ZN(n7010) );
  CKND2D0BWP U9087 ( .A1(n5865), .A2(cycles[3]), .ZN(n7011) );
  CKND0BWP U9088 ( .I(N3436), .ZN(n7009) );
  OAI22D0BWP U9089 ( .A1(n7008), .A2(n7012), .B1(n2522), .B2(n7013), .ZN(N4068) );
  CKXOR2D0BWP U9090 ( .A1(n5865), .A2(n5879), .Z(n7013) );
  CKND0BWP U9091 ( .I(cycles[3]), .ZN(n5879) );
  NR2D0BWP U9092 ( .A1(n5874), .A2(n5869), .ZN(n5865) );
  CKND0BWP U9093 ( .I(cycles[2]), .ZN(n5869) );
  CKND0BWP U9094 ( .I(N3435), .ZN(n7012) );
  OAI22D0BWP U9095 ( .A1(n7008), .A2(n7014), .B1(n2522), .B2(n7015), .ZN(N4067) );
  CKXOR2D0BWP U9096 ( .A1(cycles[2]), .A2(n5874), .Z(n7015) );
  CKND2D0BWP U9097 ( .A1(cycles[1]), .A2(cycles[0]), .ZN(n5874) );
  OAI22D0BWP U9098 ( .A1(n7008), .A2(n7016), .B1(n2522), .B2(n7017), .ZN(N4066) );
  AOI21D0BWP U9099 ( .A1(cycles[1]), .A2(n5866), .B(n5856), .ZN(n7017) );
  NR2D0BWP U9100 ( .A1(n5866), .A2(cycles[1]), .ZN(n5856) );
  OAI22D0BWP U9101 ( .A1(cycles[0]), .A2(n2522), .B1(n7008), .B2(n7018), .ZN(
        N4065) );
  OAI211D0BWP U9102 ( .A1(n2522), .A2(n6168), .B(n3262), .C(n6157), .ZN(N4064)
         );
  AOI21D0BWP U9103 ( .A1(n7019), .A2(N4105), .B(n7020), .ZN(n6157) );
  CKND2D0BWP U9104 ( .A1(n6205), .A2(n6197), .ZN(N4105) );
  OAI22D0BWP U9105 ( .A1(n6180), .A2(n7021), .B1(n6186), .B2(n7022), .ZN(N4063) );
  OAI22D0BWP U9106 ( .A1(n6180), .A2(n7023), .B1(n6187), .B2(n7022), .ZN(N4062) );
  OAI22D0BWP U9107 ( .A1(n6180), .A2(n7024), .B1(n6188), .B2(n7022), .ZN(N4061) );
  OAI22D0BWP U9108 ( .A1(n6180), .A2(n7025), .B1(n6189), .B2(n7022), .ZN(N4060) );
  OAI22D0BWP U9109 ( .A1(n6180), .A2(n7026), .B1(n6190), .B2(n7022), .ZN(N4059) );
  OAI22D0BWP U9110 ( .A1(n6180), .A2(n7027), .B1(n6191), .B2(n7022), .ZN(N4058) );
  OAI22D0BWP U9111 ( .A1(n6180), .A2(n7028), .B1(n5989), .B2(n7022), .ZN(N4057) );
  OAI22D0BWP U9112 ( .A1(n6180), .A2(n7029), .B1(n5990), .B2(n7022), .ZN(N4056) );
  OAI22D0BWP U9113 ( .A1(n6180), .A2(n7030), .B1(n5991), .B2(n7022), .ZN(N4055) );
  OAI22D0BWP U9114 ( .A1(n6180), .A2(n7031), .B1(n5992), .B2(n7022), .ZN(N4054) );
  OAI22D0BWP U9115 ( .A1(n6180), .A2(n7032), .B1(n5993), .B2(n7022), .ZN(N4053) );
  OAI22D0BWP U9116 ( .A1(n7033), .A2(n6180), .B1(n5994), .B2(n7022), .ZN(N4052) );
  OAI22D0BWP U9117 ( .A1(n7034), .A2(n6180), .B1(n5995), .B2(n7022), .ZN(N4051) );
  OAI22D0BWP U9118 ( .A1(n7035), .A2(n6180), .B1(n5996), .B2(n7022), .ZN(N4050) );
  OAI22D0BWP U9119 ( .A1(n7036), .A2(n6180), .B1(n5997), .B2(n7022), .ZN(N4049) );
  OAI22D0BWP U9120 ( .A1(n7037), .A2(n6180), .B1(n5998), .B2(n7022), .ZN(N4048) );
  OAI211D0BWP U9121 ( .A1(n7039), .A2(n7040), .B(n3266), .C(n7436), .ZN(N4047)
         );
  CKND0BWP U9122 ( .I(Reset), .ZN(n7436) );
  CKND2D0BWP U9123 ( .A1(n7038), .A2(n5544), .ZN(n7040) );
  OAI22D0BWP U9124 ( .A1(n6180), .A2(n3392), .B1(n6171), .B2(n7021), .ZN(N4044) );
  CKND0BWP U9125 ( .I(N222), .ZN(n7021) );
  OAI22D0BWP U9126 ( .A1(n6180), .A2(n3393), .B1(n6171), .B2(n7023), .ZN(N4043) );
  CKND0BWP U9127 ( .I(N221), .ZN(n7023) );
  OAI22D0BWP U9128 ( .A1(n6180), .A2(n3394), .B1(n6171), .B2(n7024), .ZN(N4042) );
  CKND0BWP U9129 ( .I(N220), .ZN(n7024) );
  OAI22D0BWP U9130 ( .A1(n6180), .A2(n3395), .B1(n6171), .B2(n7025), .ZN(N4041) );
  CKND0BWP U9131 ( .I(N219), .ZN(n7025) );
  OAI22D0BWP U9132 ( .A1(n6180), .A2(n3396), .B1(n6171), .B2(n7026), .ZN(N4040) );
  CKND0BWP U9133 ( .I(N218), .ZN(n7026) );
  OAI22D0BWP U9134 ( .A1(n6180), .A2(n3397), .B1(n6171), .B2(n7027), .ZN(N4039) );
  CKND0BWP U9135 ( .I(N217), .ZN(n7027) );
  OAI22D0BWP U9136 ( .A1(n6180), .A2(n3398), .B1(n6171), .B2(n7028), .ZN(N4038) );
  CKND0BWP U9137 ( .I(N216), .ZN(n7028) );
  OAI22D0BWP U9138 ( .A1(n6180), .A2(n3399), .B1(n6171), .B2(n7029), .ZN(N4037) );
  CKND0BWP U9139 ( .I(N215), .ZN(n7029) );
  OAI22D0BWP U9140 ( .A1(n6180), .A2(n3400), .B1(n6171), .B2(n7030), .ZN(N4036) );
  CKND0BWP U9141 ( .I(N214), .ZN(n7030) );
  OAI22D0BWP U9142 ( .A1(n6180), .A2(n3401), .B1(n6171), .B2(n7031), .ZN(N4035) );
  CKND0BWP U9143 ( .I(N213), .ZN(n7031) );
  OAI22D0BWP U9144 ( .A1(n6180), .A2(n3402), .B1(n6171), .B2(n7032), .ZN(N4034) );
  CKND0BWP U9145 ( .I(N212), .ZN(n7032) );
  OAI22D0BWP U9146 ( .A1(n6180), .A2(n3420), .B1(n6171), .B2(n7033), .ZN(N4033) );
  OAI22D0BWP U9147 ( .A1(n6180), .A2(n3421), .B1(n6171), .B2(n7034), .ZN(N4032) );
  OAI22D0BWP U9148 ( .A1(n6180), .A2(n3422), .B1(n6171), .B2(n7035), .ZN(N4031) );
  OAI22D0BWP U9149 ( .A1(n6180), .A2(n3423), .B1(n6171), .B2(n7036), .ZN(N4030) );
  OAI22D0BWP U9150 ( .A1(n6180), .A2(n3424), .B1(n6171), .B2(n7037), .ZN(N4029) );
  CKND2D0BWP U9151 ( .A1(n6171), .A2(n3266), .ZN(N4028) );
  CKND0BWP U9152 ( .I(n5574), .ZN(WR) );
  MUX2ND0BWP U9153 ( .I0(n6186), .I1(n7042), .S(n7043), .ZN(N3768) );
  CKMUX2D0BWP U9154 ( .I0(scalarToLoad[14]), .I1(result[14]), .S(n5986), .Z(
        N3767) );
  MUX2ND0BWP U9155 ( .I0(n6188), .I1(n7044), .S(n7043), .ZN(N3766) );
  MUX2ND0BWP U9156 ( .I0(n6189), .I1(n7045), .S(n7043), .ZN(N3765) );
  MUX2ND0BWP U9157 ( .I0(n6190), .I1(n7046), .S(n7043), .ZN(N3764) );
  MUX2ND0BWP U9158 ( .I0(n6191), .I1(n7047), .S(n7043), .ZN(N3763) );
  MUX2ND0BWP U9159 ( .I0(n5989), .I1(n3390), .S(n7043), .ZN(N3762) );
  MUX2ND0BWP U9160 ( .I0(n5990), .I1(n3391), .S(n7043), .ZN(N3761) );
  MUX2ND0BWP U9161 ( .I0(n5991), .I1(n3382), .S(n7043), .ZN(N3760) );
  MUX2ND0BWP U9162 ( .I0(n5992), .I1(n3383), .S(n7043), .ZN(N3759) );
  MUX2ND0BWP U9163 ( .I0(n5993), .I1(n3384), .S(n7043), .ZN(N3758) );
  MUX2ND0BWP U9164 ( .I0(n5994), .I1(n3385), .S(n7043), .ZN(N3757) );
  MUX2ND0BWP U9165 ( .I0(n5995), .I1(n3386), .S(n7043), .ZN(N3756) );
  MUX2ND0BWP U9166 ( .I0(n5996), .I1(n3387), .S(n7043), .ZN(N3755) );
  MUX2ND0BWP U9167 ( .I0(n5997), .I1(n3388), .S(n7043), .ZN(N3754) );
  MUX2ND0BWP U9168 ( .I0(n5998), .I1(n3389), .S(n7043), .ZN(N3753) );
  INR3D0BWP U9169 ( .A1(n7048), .B1(n7049), .B2(n6215), .ZN(N2626) );
  OAI22D0BWP U9170 ( .A1(n7050), .A2(n6186), .B1(n7051), .B2(n7042), .ZN(N1762) );
  CKND0BWP U9171 ( .I(scalarToLoad[15]), .ZN(n7042) );
  AOI22D0BWP U9172 ( .A1(n7052), .A2(n5987), .B1(n7053), .B2(n6196), .ZN(n7051) );
  CKND0BWP U9173 ( .I(result[15]), .ZN(n6186) );
  NR2D0BWP U9174 ( .A1(n7054), .A2(n6210), .ZN(n7050) );
  AOI21D0BWP U9175 ( .A1(n5987), .A2(n7055), .B(n7053), .ZN(n7054) );
  CKND0BWP U9176 ( .I(n7056), .ZN(n7053) );
  OAI211D0BWP U9177 ( .A1(n6160), .A2(n7057), .B(n7058), .C(n7059), .ZN(N1761)
         );
  AOI22D0BWP U9178 ( .A1(n7060), .A2(N3436), .B1(n6210), .B2(result[14]), .ZN(
        n7059) );
  MUX2ND0BWP U9179 ( .I0(n7061), .I1(N1565), .S(n7062), .ZN(n6160) );
  OAI211D0BWP U9180 ( .A1(n6161), .A2(n7057), .B(n7058), .C(n7063), .ZN(N1760)
         );
  AOI22D0BWP U9181 ( .A1(n7060), .A2(N3435), .B1(n6210), .B2(result[13]), .ZN(
        n7063) );
  MUX2ND0BWP U9182 ( .I0(n7064), .I1(n7065), .S(n7066), .ZN(n6161) );
  OAI211D0BWP U9183 ( .A1(n6162), .A2(n7057), .B(n7058), .C(n7067), .ZN(N1759)
         );
  AOI22D0BWP U9184 ( .A1(n7060), .A2(N3434), .B1(n6210), .B2(result[12]), .ZN(
        n7067) );
  MUX2ND0BWP U9185 ( .I0(n7068), .I1(N1563), .S(n7062), .ZN(n6162) );
  OAI211D0BWP U9186 ( .A1(n6163), .A2(n7057), .B(n7058), .C(n7069), .ZN(N1758)
         );
  AOI22D0BWP U9187 ( .A1(n7060), .A2(N3433), .B1(n6210), .B2(result[11]), .ZN(
        n7069) );
  MUX2ND0BWP U9188 ( .I0(n7070), .I1(N1562), .S(n7062), .ZN(n6163) );
  OAI211D0BWP U9189 ( .A1(n6164), .A2(n7057), .B(n7058), .C(n7071), .ZN(N1757)
         );
  AOI22D0BWP U9190 ( .A1(n7060), .A2(N3432), .B1(n6210), .B2(result[10]), .ZN(
        n7071) );
  OA21D0BWP U9191 ( .A1(n6166), .A2(n6167), .B(n7052), .Z(n7060) );
  CKND2D0BWP U9192 ( .A1(n6196), .A2(n7072), .ZN(n7058) );
  CKND2D0BWP U9193 ( .A1(n7073), .A2(n7052), .ZN(n7057) );
  MUX2ND0BWP U9194 ( .I0(n7074), .I1(N1561), .S(n7062), .ZN(n6164) );
  OAI22D0BWP U9195 ( .A1(n5989), .A2(n6196), .B1(n7075), .B2(n7076), .ZN(N1756) );
  AOI222D0BWP U9196 ( .A1(n7077), .A2(n6166), .B1(N1691), .B2(n6167), .C1(
        n7449), .C2(n7073), .ZN(n7075) );
  CKND0BWP U9197 ( .I(result[9]), .ZN(n5989) );
  OAI22D0BWP U9198 ( .A1(n5990), .A2(n6196), .B1(n7078), .B2(n7076), .ZN(N1755) );
  AOI222D0BWP U9199 ( .A1(n7449), .A2(n6166), .B1(N1690), .B2(n6167), .C1(
        n7073), .C2(N1610), .ZN(n7078) );
  CKND0BWP U9200 ( .I(result[8]), .ZN(n5990) );
  OAI22D0BWP U9201 ( .A1(n5991), .A2(n6196), .B1(n7079), .B2(n7076), .ZN(N1754) );
  AOI222D0BWP U9202 ( .A1(n6166), .A2(N1610), .B1(N1689), .B2(n6167), .C1(
        n7448), .C2(n7073), .ZN(n7079) );
  CKND0BWP U9203 ( .I(result[7]), .ZN(n5991) );
  OAI22D0BWP U9204 ( .A1(n5992), .A2(n6196), .B1(n7080), .B2(n7076), .ZN(N1753) );
  AOI222D0BWP U9205 ( .A1(n7448), .A2(n6166), .B1(N1688), .B2(n6167), .C1(
        n7447), .C2(n7073), .ZN(n7080) );
  CKND0BWP U9206 ( .I(result[6]), .ZN(n5992) );
  OAI22D0BWP U9207 ( .A1(n5993), .A2(n6196), .B1(n7081), .B2(n7076), .ZN(N1752) );
  AOI222D0BWP U9208 ( .A1(n7447), .A2(n6166), .B1(N1687), .B2(n6167), .C1(
        n7446), .C2(n7073), .ZN(n7081) );
  CKND0BWP U9209 ( .I(result[5]), .ZN(n5993) );
  OAI22D0BWP U9210 ( .A1(n5994), .A2(n6196), .B1(n7082), .B2(n7076), .ZN(N1751) );
  AOI222D0BWP U9211 ( .A1(n7446), .A2(n6166), .B1(N1686), .B2(n6167), .C1(
        n7445), .C2(n7073), .ZN(n7082) );
  CKND0BWP U9212 ( .I(result[4]), .ZN(n5994) );
  OAI22D0BWP U9213 ( .A1(n5995), .A2(n6196), .B1(n7083), .B2(n7076), .ZN(N1750) );
  AOI222D0BWP U9214 ( .A1(n7445), .A2(n6166), .B1(N1685), .B2(n6167), .C1(
        n7444), .C2(n7073), .ZN(n7083) );
  CKND0BWP U9215 ( .I(result[3]), .ZN(n5995) );
  OAI22D0BWP U9216 ( .A1(n5996), .A2(n6196), .B1(n7084), .B2(n7076), .ZN(N1749) );
  AOI222D0BWP U9217 ( .A1(n7444), .A2(n6166), .B1(N1684), .B2(n6167), .C1(
        n7443), .C2(n7073), .ZN(n7084) );
  CKND0BWP U9218 ( .I(result[2]), .ZN(n5996) );
  OAI22D0BWP U9219 ( .A1(n5997), .A2(n6196), .B1(n7085), .B2(n7076), .ZN(N1748) );
  AOI222D0BWP U9220 ( .A1(n7443), .A2(n6166), .B1(N1683), .B2(n6167), .C1(
        n7073), .C2(n7442), .ZN(n7085) );
  CKND0BWP U9221 ( .I(n6152), .ZN(n7443) );
  CKND0BWP U9222 ( .I(result[1]), .ZN(n5997) );
  OAI22D0BWP U9223 ( .A1(n5998), .A2(n6196), .B1(n7086), .B2(n7076), .ZN(N1747) );
  IND2D0BWP U9224 ( .A1(n7072), .B1(n7052), .ZN(n7076) );
  NR2D0BWP U9225 ( .A1(n6210), .A2(n6251), .ZN(n7052) );
  CKND0BWP U9226 ( .I(n7055), .ZN(n6251) );
  CKND0BWP U9227 ( .I(n6196), .ZN(n6210) );
  ND4D0BWP U9228 ( .A1(n7055), .A2(n7087), .A3(n7056), .A4(n7088), .ZN(n7072)
         );
  AOI31D0BWP U9229 ( .A1(n7089), .A2(n7065), .A3(n7090), .B(n7091), .ZN(n7088)
         );
  NR4D0BWP U9230 ( .A1(n7092), .A2(n7018), .A3(n7014), .A4(n7016), .ZN(n7091)
         );
  CKND0BWP U9231 ( .I(N3433), .ZN(n7016) );
  CKND0BWP U9232 ( .I(N3434), .ZN(n7014) );
  CKND0BWP U9233 ( .I(N3432), .ZN(n7018) );
  ND3D0BWP U9234 ( .A1(N3436), .A2(n6166), .A3(N3435), .ZN(n7092) );
  AN2D0BWP U9235 ( .A1(n7455), .A2(n7093), .Z(n7090) );
  CKMUX2D0BWP U9236 ( .I0(n7064), .I1(N1564), .S(n7094), .Z(n7065) );
  MUX2ND0BWP U9237 ( .I0(n7095), .I1(n7096), .S(n7094), .ZN(n7089) );
  ND4D0BWP U9238 ( .A1(N1561), .A2(N1562), .A3(N1563), .A4(N1565), .ZN(n7096)
         );
  ND4D0BWP U9239 ( .A1(n7074), .A2(n7061), .A3(n7068), .A4(n7070), .ZN(n7095)
         );
  AOI222D0BWP U9240 ( .A1(n7442), .A2(n6166), .B1(N1682), .B2(n6167), .C1(
        n7073), .C2(N1602), .ZN(n7086) );
  NR2D0BWP U9241 ( .A1(n7097), .A2(n6166), .ZN(n7073) );
  INR3D0BWP U9242 ( .A1(n7098), .B1(n6166), .B2(n7077), .ZN(n6167) );
  CKND0BWP U9243 ( .I(n7097), .ZN(n7077) );
  MUX2ND0BWP U9244 ( .I0(N1537), .I1(N1557), .S(n7066), .ZN(n7097) );
  ND4D0BWP U9245 ( .A1(n6147), .A2(n6153), .A3(n7099), .A4(n6152), .ZN(n7098)
         );
  INR4D0BWP U9246 ( .A1(n7100), .B1(n7449), .B2(N1610), .B3(n7448), .ZN(n6147)
         );
  CKND0BWP U9247 ( .I(n6155), .ZN(n6166) );
  CKND2D0BWP U9248 ( .A1(N1558), .A2(n7066), .ZN(n6155) );
  ND3D0BWP U9249 ( .A1(n5866), .A2(n5868), .A3(n5857), .ZN(n6196) );
  INR2D0BWP U9250 ( .A1(n5863), .B1(cycles[2]), .ZN(n5857) );
  NR2D0BWP U9251 ( .A1(cycles[4]), .A2(cycles[3]), .ZN(n5863) );
  CKND0BWP U9252 ( .I(cycles[1]), .ZN(n5868) );
  CKND0BWP U9253 ( .I(result[0]), .ZN(n5998) );
  AOI21D0BWP U9254 ( .A1(n7102), .A2(n7103), .B(n7448), .ZN(n7101) );
  OAI21D0BWP U9255 ( .A1(n7104), .A2(n7445), .B(n7105), .ZN(n7103) );
  AOI21D0BWP U9256 ( .A1(n7442), .A2(n6152), .B(n7444), .ZN(n7104) );
  MUX2ND0BWP U9257 ( .I0(N1529), .I1(N1549), .S(n7066), .ZN(n6152) );
  CKND0BWP U9258 ( .I(n6153), .ZN(n7442) );
  MUX2ND0BWP U9259 ( .I0(N1528), .I1(N1548), .S(n7066), .ZN(n6153) );
  NR4D0BWP U9260 ( .A1(n7447), .A2(n7446), .A3(n7445), .A4(n7444), .ZN(n7100)
         );
  CKMUX2D0BWP U9261 ( .I0(N1530), .I1(N1550), .S(n7066), .Z(n7444) );
  CKND0BWP U9262 ( .I(n6151), .ZN(n7445) );
  MUX2ND0BWP U9263 ( .I0(N1531), .I1(N1551), .S(n7066), .ZN(n6151) );
  CKND0BWP U9264 ( .I(n7105), .ZN(n7446) );
  MUX2ND0BWP U9265 ( .I0(N1532), .I1(N1552), .S(n7066), .ZN(n7105) );
  CKND0BWP U9266 ( .I(n7102), .ZN(n7447) );
  MUX2ND0BWP U9267 ( .I0(N1533), .I1(N1553), .S(n7066), .ZN(n7102) );
  CKMUX2D0BWP U9268 ( .I0(N1534), .I1(N1554), .S(n7066), .Z(n7448) );
  CKND0BWP U9269 ( .I(n6149), .ZN(n7449) );
  MUX2ND0BWP U9270 ( .I0(N1536), .I1(N1556), .S(n7066), .ZN(n6149) );
  CKMUX2D0BWP U9271 ( .I0(N1535), .I1(N1555), .S(n7066), .Z(N1610) );
  CKND0BWP U9272 ( .I(n7099), .ZN(N1602) );
  MUX2ND0BWP U9273 ( .I0(N1527), .I1(N1547), .S(n7066), .ZN(n7099) );
  CKMUX2D0BWP U9274 ( .I0(n7455), .I1(N1546), .S(n7066), .Z(N1601) );
  CKMUX2D0BWP U9275 ( .I0(n7454), .I1(N1545), .S(n7066), .Z(N1600) );
  XOR3D0BWP U9276 ( .A1(n6204), .A2(n7049), .A3(n7048), .Z(N1565) );
  MAOI222D0BWP U9277 ( .A(n6204), .B(n7106), .C(n7107), .ZN(n7048) );
  AOI22D0BWP U9278 ( .A1(n6215), .A2(n7108), .B1(n7109), .B2(n7110), .ZN(n7106) );
  OR2D0BWP U9279 ( .A1(n7110), .A2(n7109), .Z(n7108) );
  CKND0BWP U9280 ( .I(n7111), .ZN(n7109) );
  AOI22D0BWP U9281 ( .A1(cycles[4]), .A2(n6215), .B1(n7061), .B2(n7112), .ZN(
        n7049) );
  OAI22D0BWP U9282 ( .A1(n7113), .A2(n7033), .B1(n6183), .B2(n7114), .ZN(n7061) );
  MUX2ND0BWP U9283 ( .I0(scalarToLoad[14]), .I1(result[14]), .S(n5988), .ZN(
        n6183) );
  XNR3D0BWP U9284 ( .A1(n6215), .A2(n7107), .A3(n7115), .ZN(N1564) );
  MAOI222D0BWP U9285 ( .A(n6204), .B(n7116), .C(n7111), .ZN(n7115) );
  MAOI22D0BWP U9286 ( .A1(n6215), .A2(n7117), .B1(n7118), .B2(N1561), .ZN(
        n7116) );
  CKND2D0BWP U9287 ( .A1(N1561), .A2(n7118), .ZN(n7117) );
  AOI22D0BWP U9288 ( .A1(cycles[3]), .A2(n6215), .B1(n7064), .B2(n7112), .ZN(
        n7107) );
  OAI22D0BWP U9289 ( .A1(n7113), .A2(n7034), .B1(n7114), .B2(n6184), .ZN(n7064) );
  MUX2ND0BWP U9290 ( .I0(scalarToLoad[13]), .I1(result[13]), .S(n5988), .ZN(
        n6184) );
  MAOI222D0BWP U9291 ( .A(n6204), .B(N1561), .C(n7118), .ZN(n7110) );
  AOI22D0BWP U9292 ( .A1(n7112), .A2(n7068), .B1(n6215), .B2(cycles[2]), .ZN(
        n7111) );
  OAI22D0BWP U9293 ( .A1(n7113), .A2(n7035), .B1(n7114), .B2(n6185), .ZN(n7068) );
  MUX2ND0BWP U9294 ( .I0(scalarToLoad[12]), .I1(result[12]), .S(n5988), .ZN(
        n6185) );
  AOI22D0BWP U9295 ( .A1(cycles[1]), .A2(n6215), .B1(n7070), .B2(n7112), .ZN(
        n7118) );
  OAI22D0BWP U9296 ( .A1(n7113), .A2(n7036), .B1(n7114), .B2(n6192), .ZN(n7070) );
  MUX2ND0BWP U9297 ( .I0(scalarToLoad[11]), .I1(result[11]), .S(n5988), .ZN(
        n6192) );
  CKND0BWP U9298 ( .I(N208), .ZN(n7036) );
  CKND0BWP U9299 ( .I(n6204), .ZN(n6215) );
  CKND2D0BWP U9300 ( .A1(n7041), .A2(n5988), .ZN(n6204) );
  AN2D0BWP U9301 ( .A1(n7062), .A2(n6195), .Z(n7112) );
  AN2D0BWP U9302 ( .A1(n7094), .A2(n7066), .Z(n7062) );
  AN3D0BWP U9303 ( .A1(n7087), .A2(n7455), .A3(n7093), .Z(n7066) );
  ND4D0BWP U9304 ( .A1(n7119), .A2(n7120), .A3(n7121), .A4(n7122), .ZN(n7093)
         );
  NR4D0BWP U9305 ( .A1(N1266), .A2(N1265), .A3(N1264), .A4(N1263), .ZN(n7122)
         );
  NR4D0BWP U9306 ( .A1(N1262), .A2(N1261), .A3(N1260), .A4(N1259), .ZN(n7121)
         );
  NR4D0BWP U9307 ( .A1(N1258), .A2(N1257), .A3(N1256), .A4(N1255), .ZN(n7120)
         );
  NR3D0BWP U9308 ( .A1(n7123), .A2(n7454), .A3(N1527), .ZN(n7119) );
  AO222D0BWP U9309 ( .A1(N1407), .A2(n7124), .B1(N1488), .B2(n6194), .C1(N1408), .C2(N1280), .Z(n7454) );
  MUX2ND0BWP U9310 ( .I0(n7125), .I1(n7126), .S(N1280), .ZN(n7123) );
  AO222D0BWP U9311 ( .A1(N1409), .A2(N1280), .B1(N1489), .B2(n6194), .C1(N1408), .C2(n7124), .Z(n7455) );
  ND4D0BWP U9312 ( .A1(N207), .A2(N1280), .A3(N208), .A4(n7127), .ZN(n7087) );
  NR3D0BWP U9313 ( .A1(n7033), .A2(n7035), .A3(n7034), .ZN(n7127) );
  CKND0BWP U9314 ( .I(N210), .ZN(n7034) );
  CKND0BWP U9315 ( .I(N209), .ZN(n7035) );
  CKND0BWP U9316 ( .I(N211), .ZN(n7033) );
  IINR4D0BWP U9317 ( .A1(n7128), .A2(n7129), .B1(N1547), .B2(N1548), .ZN(n7094) );
  NR4D0BWP U9318 ( .A1(n7130), .A2(N1554), .A3(N1556), .A4(N1555), .ZN(n7129)
         );
  OR2D0BWP U9319 ( .A1(N1552), .A2(N1553), .Z(n7130) );
  NR3D0BWP U9320 ( .A1(N1549), .A2(N1551), .A3(N1550), .ZN(n7128) );
  OAI22D0BWP U9321 ( .A1(n7113), .A2(n7037), .B1(n6193), .B2(n7114), .ZN(n7074) );
  MUX2ND0BWP U9322 ( .I0(result[10]), .I1(scalarToLoad[10]), .S(n5987), .ZN(
        n6193) );
  CKND2D0BWP U9323 ( .A1(n7131), .A2(n7132), .ZN(n5988) );
  AO21D0BWP U9324 ( .A1(scalarToLoad[14]), .A2(n6195), .B(n7133), .Z(n7132) );
  OAI32D0BWP U9325 ( .A1(n7134), .A2(n7135), .A3(n7136), .B1(n7137), .B2(n7138), .ZN(n7131) );
  AOI22D0BWP U9326 ( .A1(n7139), .A2(scalarToLoad[13]), .B1(n7133), .B2(
        scalarToLoad[14]), .ZN(n7137) );
  AOI22D0BWP U9327 ( .A1(n7041), .A2(cycles[4]), .B1(result[14]), .B2(n6195), 
        .ZN(n7133) );
  AOI21D0BWP U9328 ( .A1(n6195), .A2(scalarToLoad[13]), .B(n7139), .ZN(n7136)
         );
  AOI22D0BWP U9329 ( .A1(cycles[3]), .A2(n7041), .B1(result[13]), .B2(n6195), 
        .ZN(n7139) );
  AOI22D0BWP U9330 ( .A1(n6195), .A2(scalarToLoad[12]), .B1(n7140), .B2(n7141), 
        .ZN(n7135) );
  NR2D0BWP U9331 ( .A1(n7140), .A2(n7141), .ZN(n7134) );
  OA32D0BWP U9332 ( .A1(n7142), .A2(n6191), .A3(n7138), .B1(n7143), .B2(n7144), 
        .Z(n7141) );
  AO21D0BWP U9333 ( .A1(n7144), .A2(n7143), .B(scalarToLoad[10]), .Z(n7142) );
  NR2D0BWP U9334 ( .A1(n7138), .A2(n7046), .ZN(n7143) );
  AOI22D0BWP U9335 ( .A1(cycles[1]), .A2(n7041), .B1(result[11]), .B2(n6195), 
        .ZN(n7144) );
  AOI22D0BWP U9336 ( .A1(cycles[2]), .A2(n7041), .B1(result[12]), .B2(n6195), 
        .ZN(n7140) );
  CKND0BWP U9337 ( .I(n7138), .ZN(n6195) );
  ND3D0BWP U9338 ( .A1(n7055), .A2(n6466), .A3(n7056), .ZN(n7138) );
  ND4D0BWP U9339 ( .A1(scalarToLoad[14]), .A2(scalarToLoad[13]), .A3(n7145), 
        .A4(scalarToLoad[12]), .ZN(n7056) );
  NR2D0BWP U9340 ( .A1(n7047), .A2(n7046), .ZN(n7145) );
  ND4D0BWP U9341 ( .A1(result[14]), .A2(result[13]), .A3(n7146), .A4(
        result[12]), .ZN(n7055) );
  NR2D0BWP U9342 ( .A1(n6191), .A2(n6190), .ZN(n7146) );
  CKND0BWP U9343 ( .I(N207), .ZN(n7037) );
  NR2D0BWP U9344 ( .A1(n6194), .A2(N1280), .ZN(n7113) );
  AO211D0BWP U9345 ( .A1(N1500), .A2(n6194), .B(N1419), .C(N1280), .Z(N1537)
         );
  AO222D0BWP U9346 ( .A1(N1418), .A2(n7124), .B1(N1499), .B2(n6194), .C1(N1419), .C2(N1280), .Z(N1536) );
  AO222D0BWP U9347 ( .A1(N1417), .A2(n7124), .B1(N1498), .B2(n6194), .C1(N1418), .C2(N1280), .Z(N1535) );
  AO222D0BWP U9348 ( .A1(N1416), .A2(n7124), .B1(N1497), .B2(n6194), .C1(N1417), .C2(N1280), .Z(N1534) );
  AO222D0BWP U9349 ( .A1(N1415), .A2(n7124), .B1(N1496), .B2(n6194), .C1(N1416), .C2(N1280), .Z(N1533) );
  AO222D0BWP U9350 ( .A1(N1414), .A2(n7124), .B1(N1495), .B2(n6194), .C1(N1415), .C2(N1280), .Z(N1532) );
  AO222D0BWP U9351 ( .A1(N1413), .A2(n7124), .B1(N1494), .B2(n6194), .C1(N1414), .C2(N1280), .Z(N1531) );
  AO222D0BWP U9352 ( .A1(N1412), .A2(n7124), .B1(N1493), .B2(n6194), .C1(N1413), .C2(N1280), .Z(N1530) );
  AO222D0BWP U9353 ( .A1(N1411), .A2(n7124), .B1(N1492), .B2(n6194), .C1(N1412), .C2(N1280), .Z(N1529) );
  AO222D0BWP U9354 ( .A1(N1410), .A2(n7124), .B1(N1491), .B2(n6194), .C1(N1411), .C2(N1280), .Z(N1528) );
  AO222D0BWP U9355 ( .A1(N1409), .A2(n7124), .B1(N1490), .B2(n6194), .C1(N1410), .C2(N1280), .Z(N1527) );
  INR3D0BWP U9356 ( .A1(n7147), .B1(N1419), .B2(N1280), .ZN(n6194) );
  CKND2D0BWP U9357 ( .A1(n7147), .A2(n7114), .ZN(n7124) );
  CKND2D0BWP U9358 ( .A1(N1419), .A2(n6179), .ZN(n7114) );
  CKND0BWP U9359 ( .I(N1280), .ZN(n6179) );
  ND4D0BWP U9360 ( .A1(n7148), .A2(n7149), .A3(n7150), .A4(n6177), .ZN(n7147)
         );
  NR2D0BWP U9361 ( .A1(N1418), .A2(N1280), .ZN(n7150) );
  MUX2ND0BWP U9362 ( .I0(n7151), .I1(n7126), .S(N1280), .ZN(N1524) );
  CKND0BWP U9363 ( .I(N1407), .ZN(n7126) );
  MUX2ND0BWP U9364 ( .I0(n7152), .I1(n7151), .S(N1280), .ZN(N1523) );
  CKND0BWP U9365 ( .I(N1266), .ZN(n7151) );
  MUX2ND0BWP U9366 ( .I0(n7153), .I1(n7152), .S(N1280), .ZN(N1522) );
  CKND0BWP U9367 ( .I(N1265), .ZN(n7152) );
  MUX2ND0BWP U9368 ( .I0(n7154), .I1(n7153), .S(N1280), .ZN(N1521) );
  CKND0BWP U9369 ( .I(N1264), .ZN(n7153) );
  MUX2ND0BWP U9370 ( .I0(n7155), .I1(n7154), .S(N1280), .ZN(N1520) );
  CKND0BWP U9371 ( .I(N1263), .ZN(n7154) );
  MUX2ND0BWP U9372 ( .I0(n5561), .I1(n7155), .S(N1280), .ZN(N1519) );
  CKND0BWP U9373 ( .I(N1262), .ZN(n7155) );
  CKND0BWP U9374 ( .I(N1261), .ZN(n5561) );
  MUX2ND0BWP U9375 ( .I0(n7156), .I1(n5557), .S(N1280), .ZN(N1514) );
  CKND0BWP U9376 ( .I(N1257), .ZN(n5557) );
  MUX2ND0BWP U9377 ( .I0(n7157), .I1(n7156), .S(N1280), .ZN(N1513) );
  CKND0BWP U9378 ( .I(N1256), .ZN(n7156) );
  MUX2ND0BWP U9379 ( .I0(n7125), .I1(n7157), .S(N1280), .ZN(N1512) );
  CKND0BWP U9380 ( .I(N1255), .ZN(n7157) );
  CKND0BWP U9381 ( .I(N1254), .ZN(n7125) );
  AOI21D0BWP U9382 ( .A1(n7159), .A2(n7160), .B(N1416), .ZN(n7158) );
  CKND0BWP U9383 ( .I(N1415), .ZN(n7160) );
  OAI21D0BWP U9384 ( .A1(N1413), .A2(n7161), .B(n7162), .ZN(n7159) );
  CKND0BWP U9385 ( .I(N1414), .ZN(n7162) );
  AOI21D0BWP U9386 ( .A1(N1410), .A2(n7163), .B(N1412), .ZN(n7161) );
  CKND0BWP U9387 ( .I(N1411), .ZN(n7163) );
  CKND0BWP U9388 ( .I(n6173), .ZN(N1457) );
  IND4D0BWP U9389 ( .A1(n7149), .B1(n7148), .B2(n6177), .B3(n6174), .ZN(n6173)
         );
  CKND0BWP U9390 ( .I(N1418), .ZN(n6174) );
  NR2D0BWP U9391 ( .A1(N1416), .A2(N1417), .ZN(n6177) );
  NR4D0BWP U9392 ( .A1(N1412), .A2(N1413), .A3(N1414), .A4(N1415), .ZN(n7148)
         );
  NR3D0BWP U9393 ( .A1(N1410), .A2(N1411), .A3(N1409), .ZN(n7149) );
  NR2D0BWP U9394 ( .A1(Reset), .A2(n7164), .ZN(N140) );
  AOI22D0BWP U9395 ( .A1(n7165), .A2(n7019), .B1(n3368), .B2(n6199), .ZN(n7164) );
  CKND2D0BWP U9396 ( .A1(n2522), .A2(n6169), .ZN(n7165) );
  AOI31D0BWP U9397 ( .A1(n7166), .A2(n6977), .A3(n6170), .B(Reset), .ZN(N139)
         );
  INR2D0BWP U9398 ( .A1(n7167), .B1(n7020), .ZN(n6170) );
  OAI21D0BWP U9399 ( .A1(n7041), .A2(n6209), .B(n7019), .ZN(n7167) );
  CKND2D0BWP U9400 ( .A1(n3368), .A2(n6470), .ZN(n6977) );
  OAI21D0BWP U9401 ( .A1(n7168), .A2(n6200), .B(n3368), .ZN(n7166) );
  IND2D0BWP U9402 ( .A1(n5549), .B1(n6472), .ZN(n6200) );
  AOI31D0BWP U9403 ( .A1(n6993), .A2(n3262), .A3(n7169), .B(Reset), .ZN(N138)
         );
  AOI32D0BWP U9404 ( .A1(n3368), .A2(n5538), .A3(n7170), .B1(n6168), .B2(n7171), .ZN(n7169) );
  CKND2D0BWP U9405 ( .A1(n7172), .A2(n6169), .ZN(n7171) );
  NR2D0BWP U9406 ( .A1(n6199), .A2(n5549), .ZN(n7170) );
  CKND0BWP U9407 ( .I(n7168), .ZN(n5538) );
  NR2D0BWP U9408 ( .A1(n6396), .A2(n6198), .ZN(n7168) );
  AN2D0BWP U9409 ( .A1(n7173), .A2(n5854), .Z(n6396) );
  CKND2D0BWP U9410 ( .A1(n7174), .A2(code[0]), .ZN(n5854) );
  ND3D0BWP U9411 ( .A1(state[0]), .A2(n7039), .A3(n7175), .ZN(n3262) );
  OAI21D0BWP U9412 ( .A1(Reset), .A2(n7176), .B(n6180), .ZN(N137) );
  ND3D0BWP U9413 ( .A1(n5544), .A2(n7039), .A3(n7175), .ZN(n3266) );
  INR4D0BWP U9414 ( .A1(n6205), .B1(n7020), .B2(n7177), .B3(n7178), .ZN(n7176)
         );
  NR2D0BWP U9415 ( .A1(n7172), .A2(n7019), .ZN(n7178) );
  NR2D0BWP U9416 ( .A1(n6466), .A2(n7041), .ZN(n7172) );
  CKND0BWP U9417 ( .I(n6197), .ZN(n7041) );
  ND3D0BWP U9418 ( .A1(n7175), .A2(n5544), .A3(state[2]), .ZN(n6197) );
  CKND0BWP U9419 ( .I(n2522), .ZN(n6466) );
  CKND2D0BWP U9420 ( .A1(n7179), .A2(n5544), .ZN(n2522) );
  CKND0BWP U9421 ( .I(state[0]), .ZN(n5544) );
  NR4D0BWP U9422 ( .A1(n5549), .A2(n7043), .A3(n6470), .A4(n6250), .ZN(n7177)
         );
  CKND0BWP U9423 ( .I(n3368), .ZN(n6250) );
  NR2D0BWP U9424 ( .A1(n5545), .A2(state[0]), .ZN(n3368) );
  CKND2D0BWP U9425 ( .A1(n7038), .A2(n7039), .ZN(n5545) );
  CKND0BWP U9426 ( .I(state[2]), .ZN(n7039) );
  NR4D0BWP U9427 ( .A1(n6471), .A2(code[0]), .A3(code[1]), .A4(code[2]), .ZN(
        n6470) );
  CKND0BWP U9428 ( .I(n5986), .ZN(n7043) );
  CKND2D0BWP U9429 ( .A1(n6199), .A2(code[0]), .ZN(n5986) );
  NR2D0BWP U9430 ( .A1(n5574), .A2(n6168), .ZN(n7020) );
  CKND0BWP U9431 ( .I(n7019), .ZN(n6168) );
  ND4D0BWP U9432 ( .A1(n7180), .A2(n7181), .A3(n7182), .A4(n7183), .ZN(n7019)
         );
  NR2D0BWP U9433 ( .A1(n7184), .A2(n7185), .ZN(n7183) );
  CKXOR2D0BWP U9434 ( .A1(n5549), .A2(cycles[4]), .Z(n7185) );
  NR2D0BWP U9435 ( .A1(n7173), .A2(code[0]), .ZN(n5549) );
  CKXOR2D0BWP U9436 ( .A1(cycles[3]), .A2(cycles[2]), .Z(n7184) );
  CKXOR2D0BWP U9437 ( .A1(cycles[1]), .A2(n5878), .Z(n7182) );
  CKXOR2D0BWP U9438 ( .A1(n5550), .A2(n5866), .Z(n7181) );
  CKND0BWP U9439 ( .I(cycles[0]), .ZN(n5866) );
  OAI21D0BWP U9440 ( .A1(n6198), .A2(n7173), .B(n5536), .ZN(n5550) );
  AN2D0BWP U9441 ( .A1(n6472), .A2(n6406), .Z(n5536) );
  CKND0BWP U9442 ( .I(n6199), .ZN(n6406) );
  NR3D0BWP U9443 ( .A1(code[2]), .A2(code[3]), .A3(code[1]), .ZN(n6199) );
  CKND2D0BWP U9444 ( .A1(n7174), .A2(n6198), .ZN(n6472) );
  NR3D0BWP U9445 ( .A1(code[2]), .A2(code[3]), .A3(n6975), .ZN(n7174) );
  ND3D0BWP U9446 ( .A1(n6975), .A2(n6471), .A3(code[2]), .ZN(n7173) );
  CKND0BWP U9447 ( .I(code[3]), .ZN(n6471) );
  CKND0BWP U9448 ( .I(code[1]), .ZN(n6975) );
  CKND0BWP U9449 ( .I(code[0]), .ZN(n6198) );
  CKXOR2D0BWP U9450 ( .A1(cycles[0]), .A2(n5878), .Z(n7180) );
  CKND2D0BWP U9451 ( .A1(cycles[2]), .A2(cycles[3]), .ZN(n5878) );
  ND3D0BWP U9452 ( .A1(n7175), .A2(state[0]), .A3(state[2]), .ZN(n5574) );
  NR2D0BWP U9453 ( .A1(state[3]), .A2(state[1]), .ZN(n7175) );
  NR2D0BWP U9454 ( .A1(n6467), .A2(n6209), .ZN(n6205) );
  CKND0BWP U9455 ( .I(n6993), .ZN(n6209) );
  ND3D0BWP U9456 ( .A1(state[0]), .A2(n7038), .A3(state[2]), .ZN(n6993) );
  INR2D0BWP U9457 ( .A1(state[1]), .B1(state[3]), .ZN(n7038) );
  CKND0BWP U9458 ( .I(n6169), .ZN(n6467) );
  CKND2D0BWP U9459 ( .A1(n7179), .A2(state[0]), .ZN(n6169) );
  INR3D0BWP U9460 ( .A1(state[3]), .B1(state[1]), .B2(state[2]), .ZN(n7179) );
  ND4D0BWP U9461 ( .A1(n6188), .A2(n6187), .A3(n6189), .A4(n7186), .ZN(N1169)
         );
  NR2D0BWP U9462 ( .A1(result[11]), .A2(result[10]), .ZN(n7186) );
  ND4D0BWP U9463 ( .A1(n7047), .A2(n7046), .A3(n7187), .A4(n7045), .ZN(N1168)
         );
  NR2D0BWP U9464 ( .A1(scalarToLoad[14]), .A2(scalarToLoad[13]), .ZN(n7187) );
  XOR3D0BWP U9465 ( .A1(scalarToLoad[14]), .A2(n6187), .A3(n7188), .Z(N1167)
         );
  MAOI222D0BWP U9466 ( .A(n7044), .B(result[13]), .C(n7189), .ZN(n7188) );
  AOI22D0BWP U9467 ( .A1(scalarToLoad[12]), .A2(n7190), .B1(n7191), .B2(n6189), 
        .ZN(n7189) );
  OR2D0BWP U9468 ( .A1(n7191), .A2(n6189), .Z(n7190) );
  CKND0BWP U9469 ( .I(scalarToLoad[13]), .ZN(n7044) );
  CKND0BWP U9470 ( .I(result[14]), .ZN(n6187) );
  XOR3D0BWP U9471 ( .A1(scalarToLoad[13]), .A2(n6188), .A3(n7192), .Z(N1166)
         );
  MAOI222D0BWP U9472 ( .A(n7045), .B(result[12]), .C(n7193), .ZN(n7192) );
  AOI22D0BWP U9473 ( .A1(scalarToLoad[11]), .A2(n7194), .B1(n7195), .B2(n6190), 
        .ZN(n7193) );
  CKND0BWP U9474 ( .I(result[11]), .ZN(n6190) );
  IND2D0BWP U9475 ( .A1(n7195), .B1(result[11]), .ZN(n7194) );
  CKND0BWP U9476 ( .I(scalarToLoad[12]), .ZN(n7045) );
  CKND0BWP U9477 ( .I(result[13]), .ZN(n6188) );
  XOR3D0BWP U9478 ( .A1(scalarToLoad[12]), .A2(n6189), .A3(n7191), .Z(N1165)
         );
  MAOI222D0BWP U9479 ( .A(n7046), .B(result[11]), .C(n7196), .ZN(n7191) );
  NR2D0BWP U9480 ( .A1(scalarToLoad[10]), .A2(n6191), .ZN(n7196) );
  CKND0BWP U9481 ( .I(result[10]), .ZN(n6191) );
  CKND0BWP U9482 ( .I(result[12]), .ZN(n6189) );
  XOR3D0BWP U9483 ( .A1(result[11]), .A2(n7046), .A3(n7195), .Z(N1164) );
  CKND0BWP U9484 ( .I(scalarToLoad[11]), .ZN(n7046) );
  OAI21D0BWP U9485 ( .A1(result[10]), .A2(n7047), .B(n7195), .ZN(N1163) );
  CKND2D0BWP U9486 ( .A1(result[10]), .A2(n7047), .ZN(n7195) );
  CKND0BWP U9487 ( .I(scalarToLoad[10]), .ZN(n7047) );
endmodule

