module ALU ();

endmodule
