module VectorRegFile ();


CHANGES
endmodule
